VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LIBRARY artistTranslator STRING "4.2.1" ;
  LIBRARY artistVersion STRING "4.2.1" ;
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.001 ;
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER Active
  TYPE MASTERSLICE ;
  #PROPERTY LEF58_TYPE "TYPE DIFFUSION ;" ;
END Active

LAYER GO1
  TYPE MASTERSLICE ;
  #PROPERTY LEF58_TYPE "TYPE DIFFUSION ;" ;
END GO1

LAYER Gate
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  #DIRECTION VERTICAL ;
  PITCH 10 ;
  WIDTH 5 ;
  OFFSET 0 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 1 
    WIDTH 3 5 ;
  MINIMUMCUT 2 WIDTH 1.5 LENGTH 1.5 WITHIN 1 ;
  RESISTANCE RPERSQ 0.0736 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.15 ;
  EDGECAPACITANCE 0.0002 ;
  DCCURRENTDENSITY AVERAGE 2 ;
  PROPERTY LEF58_TYPE "TYPE POLYROUTING ;" ;
END Gate

LAYER Cont
  TYPE CUT ;
  SPACING 0.5 ;
  WIDTH 0.5 ;
  RESISTANCE 3.3 ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Cont

LAYER Metal1
  TYPE ROUTING ;
  #DIRECTION HORIZONTAL ;
  DIRECTION VERTICAL ;
  PITCH 10 ;
  WIDTH 5 ;
  OFFSET 5 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 1 
    WIDTH 3 5 ;
  MINIMUMCUT 2 WIDTH 1.5 FROMABOVE LENGTH 1.5 WITHIN 1 ;
  MINIMUMCUT 2 WIDTH 1.5 FROMBELOW LENGTH 1.5 WITHIN 1 ;
  RESISTANCE RPERSQ 0.0604 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.18 ;
  EDGECAPACITANCE 0.0002 ;
  DCCURRENTDENSITY AVERAGE 2 ;
END Metal1

LAYER Contact
  TYPE CUT ;
  SPACING 0.5 ;
  SPACING 1.1 LAYER Gate ;
  WIDTH 0.5 ;
  RESISTANCE 5 ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Contact

LAYER NSD
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  #DIRECTION VERTICAL ; 
  PITCH 10 ;
  WIDTH 5 ;
  OFFSET 0 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 1 
    WIDTH 3 5 ;
  MINIMUMCUT 2 WIDTH 1.5 LENGTH 1.5 WITHIN 1 ;
  RESISTANCE RPERSQ 0.0604 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.18 ;
  EDGECAPACITANCE 0.0002 ;
  DCCURRENTDENSITY AVERAGE 2 ;
END NSD

VIARULE Gate_Metal1 GENERATE DEFAULT
  LAYER Gate ;
    ENCLOSURE 1 1 ;
  LAYER Metal1 ;
    ENCLOSURE 1 1 ;
  LAYER Cont ;
    RECT -0.5 -0.5 0.5 0.5 ;
    SPACING 2 BY 2 ;
    RESISTANCE 0.040000 ;
END Gate_Metal1

VIARULE Metal1_NSD GENERATE DEFAULT
  LAYER Metal1 ;
    ENCLOSURE 1 1 ;
  LAYER NSD ;
    ENCLOSURE 1 1 ;
  LAYER Contact ;
    RECT -0.5 -0.5 0.5 0.5 ;
    SPACING 2 BY 2 ;
    RESISTANCE 0.200000 ;
END Metal1_NSD

VIA Gate_Metal1_0 DEFAULT
  VIARULE Gate_Metal1 ;
  CUTSIZE 1 1 ;
  LAYERS Gate Cont Metal1 ;
  CUTSPACING 1 1 ;
  ENCLOSURE 1 1 1 1 ;
  ROWCOL 2 2 ;
END Gate_Metal1_0

VIA Metal1_NSD_0 DEFAULT 
  VIARULE Metal1_NSD ;
  CUTSIZE 1 1 ;
  LAYERS Metal1 Contact NSD ;
  CUTSPACING 1 1 ;
  ENCLOSURE 1 1 1 1 ;
  ROWCOL 2 2 ;
END Metal1_NSD_0

NONDEFAULTRULE virtuosoDefaultSetup
  LAYER Gate
    WIDTH 5 ;
  END Gate
  LAYER Metal1
    WIDTH 5 ;
  END Metal1
  LAYER NSD
    WIDTH 5 ;
  END NSD
  USEVIARULE Gate_Metal1 ;
  USEVIARULE Metal1_NSD ;
END virtuosoDefaultSetup

NONDEFAULTRULE VLMDefaultSetup
  LAYER Gate
    WIDTH 5 ;
  END Gate
  LAYER Metal1
    WIDTH 5 ;
  END Metal1
  LAYER NSD
    WIDTH 5 ;
  END NSD
  USEVIARULE Gate_Metal1 ;
  USEVIARULE Metal1_NSD ;
END VLMDefaultSetup

SITE CoreSite
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 10 BY 280 ;
END CoreSite


MACRO MoS2And
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MoS2And 0 0 ;
  SIZE 340 BY 280 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 99 45 111 105 ;
        RECT 79 45 111 55 ;
        RECT 39 122 91 134 ;
        RECT 79 45 91 134 ;
        RECT 39 122 51 205 ;
      LAYER Metal1 ;
        RECT 40.695 196.625 48.695 215.85 ;
      LAYER NSD ;
        RECT 40.695 207.85 48.695 215.85 ;
      LAYER Cont ;
        RECT 41.195 203.125 42.195 204.125 ;
        RECT 41.195 201.125 42.195 202.125 ;
        RECT 41.195 199.125 42.195 200.125 ;
        RECT 41.195 197.125 42.195 198.125 ;
        RECT 43.195 203.125 44.195 204.125 ;
        RECT 43.195 201.125 44.195 202.125 ;
        RECT 43.195 199.125 44.195 200.125 ;
        RECT 43.195 197.125 44.195 198.125 ;
        RECT 45.195 203.125 46.195 204.125 ;
        RECT 45.195 201.125 46.195 202.125 ;
        RECT 45.195 199.125 46.195 200.125 ;
        RECT 45.195 197.125 46.195 198.125 ;
        RECT 47.195 203.125 48.195 204.125 ;
        RECT 47.195 201.125 48.195 202.125 ;
        RECT 47.195 199.125 48.195 200.125 ;
        RECT 47.195 197.125 48.195 198.125 ;
      LAYER Contact ;
        RECT 41.195 214.35 42.195 215.35 ;
        RECT 41.195 212.35 42.195 213.35 ;
        RECT 41.195 210.35 42.195 211.35 ;
        RECT 41.195 208.35 42.195 209.35 ;
        RECT 43.195 214.35 44.195 215.35 ;
        RECT 43.195 212.35 44.195 213.35 ;
        RECT 43.195 210.35 44.195 211.35 ;
        RECT 43.195 208.35 44.195 209.35 ;
        RECT 45.195 214.35 46.195 215.35 ;
        RECT 45.195 212.35 46.195 213.35 ;
        RECT 45.195 210.35 46.195 211.35 ;
        RECT 45.195 208.35 46.195 209.35 ;
        RECT 47.195 214.35 48.195 215.35 ;
        RECT 47.195 212.35 48.195 213.35 ;
        RECT 47.195 210.35 48.195 211.35 ;
        RECT 47.195 208.35 48.195 209.35 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 39 45 51 105 ;
        RECT 19 45 51 55 ;
        RECT 19 45 31 205 ;
      LAYER Metal1 ;
        RECT 31.035 33.42 39.035 54.12 ;
      LAYER NSD ;
        RECT 31.035 33.42 39.035 41.42 ;
      LAYER Cont ;
        RECT 31.535 52.62 32.535 53.62 ;
        RECT 31.535 50.62 32.535 51.62 ;
        RECT 31.535 48.62 32.535 49.62 ;
        RECT 31.535 46.62 32.535 47.62 ;
        RECT 33.535 52.62 34.535 53.62 ;
        RECT 33.535 50.62 34.535 51.62 ;
        RECT 33.535 48.62 34.535 49.62 ;
        RECT 33.535 46.62 34.535 47.62 ;
        RECT 35.535 52.62 36.535 53.62 ;
        RECT 35.535 50.62 36.535 51.62 ;
        RECT 35.535 48.62 36.535 49.62 ;
        RECT 35.535 46.62 36.535 47.62 ;
        RECT 37.535 52.62 38.535 53.62 ;
        RECT 37.535 50.62 38.535 51.62 ;
        RECT 37.535 48.62 38.535 49.62 ;
        RECT 37.535 46.62 38.535 47.62 ;
      LAYER Contact ;
        RECT 31.535 39.92 32.535 40.92 ;
        RECT 31.535 37.92 32.535 38.92 ;
        RECT 31.535 35.92 32.535 36.92 ;
        RECT 31.535 33.92 32.535 34.92 ;
        RECT 33.535 39.92 34.535 40.92 ;
        RECT 33.535 37.92 34.535 38.92 ;
        RECT 33.535 35.92 34.535 36.92 ;
        RECT 33.535 33.92 34.535 34.92 ;
        RECT 35.535 39.92 36.535 40.92 ;
        RECT 35.535 37.92 36.535 38.92 ;
        RECT 35.535 35.92 36.535 36.92 ;
        RECT 35.535 33.92 36.535 34.92 ;
        RECT 37.535 39.92 38.535 40.92 ;
        RECT 37.535 37.92 38.535 38.92 ;
        RECT 37.535 35.92 38.535 36.92 ;
        RECT 37.535 33.92 38.535 34.92 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 10 0 20 190 ;
    END
    PORT
      LAYER NSD ;
        RECT 50 0 60 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 200 0 210 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 0 340 20 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Contact ;
        RECT 313 211.225 314 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 313 213.225 314 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 313 215.225 314 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 313 217.225 314 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 313 261.65 314 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 313 263.65 314 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 313 265.65 314 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 313 267.65 314 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 311 211.225 312 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 311 213.225 312 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 311 215.225 312 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 311 217.225 312 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 311 261.65 312 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 311 263.65 312 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 311 265.65 312 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 311 267.65 312 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 309 211.225 310 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 309 213.225 310 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 309 215.225 310 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 309 217.225 310 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 309 261.65 310 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 309 263.65 310 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 309 265.65 310 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 309 267.65 310 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 307 211.225 308 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 307 213.225 308 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 307 215.225 308 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 307 217.225 308 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 307 261.65 308 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 307 263.65 308 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 307 265.65 308 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 307 267.65 308 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.465 212.915 172.465 213.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.465 214.915 172.465 215.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.465 216.915 172.465 217.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.465 218.915 172.465 219.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.465 261.91 172.465 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.465 263.91 172.465 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.465 265.91 172.465 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.465 267.91 172.465 268.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.465 212.915 170.465 213.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.465 214.915 170.465 215.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.465 216.915 170.465 217.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.465 218.915 170.465 219.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.465 261.91 170.465 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.465 263.91 170.465 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.465 265.91 170.465 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.465 267.91 170.465 268.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.465 212.915 168.465 213.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.465 214.915 168.465 215.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.465 216.915 168.465 217.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.465 218.915 168.465 219.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.465 261.91 168.465 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.465 263.91 168.465 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.465 265.91 168.465 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.465 267.91 168.465 268.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 165.465 212.915 166.465 213.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 165.465 214.915 166.465 215.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 165.465 216.915 166.465 217.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 165.465 218.915 166.465 219.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 165.465 261.91 166.465 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 165.465 263.91 166.465 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 165.465 265.91 166.465 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 165.465 267.91 166.465 268.91 ;
    END
    PORT
      LAYER NSD ;
        RECT 150 60 160 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 150 98.9 173.85 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 163.85 98.9 173.85 220.75 ;
    END
    PORT
      LAYER NSD ;
        RECT 240 60 250 105.55 ;
    END
    PORT
      LAYER NSD ;
        RECT 240 95.55 315.45 105.55 ;
    END
    PORT
      LAYER NSD ;
        RECT 305.45 95.55 315.45 219.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 260 340 280 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 164.965 212.415 172.965 269.41 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 306.5 210.725 314.5 269.15 ;
    END
  END VDD
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER NSD ;
        RECT 220 31.785 230 90 ;
    END
  END VOUT
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 70 160 80 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 110 160 120 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 150 160 160 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 70 198.1 160 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 200 160 210 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 240 160 250 208.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 280 160 290 208.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 200 198.95 290 208.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 230 340 250 ;
    END
  END VSS
  OBS
    LAYER Gate ;
      RECT 249 195 281 205 ;
      RECT 269 145 281 205 ;
      RECT 209 195 241 205 ;
      RECT 229 45 241 205 ;
      RECT 189 145 201 205 ;
      RECT 249 145 261 205 ;
      RECT 209 145 221 205 ;
      RECT 229 145 261 155 ;
      RECT 189 145 221 155 ;
      RECT 195 114.75 241 124.75 ;
      RECT 209 43.35 221 105 ;
      RECT 189 43.35 201 105 ;
      RECT 189 43.35 221 55.35 ;
      RECT 119 195 151 205 ;
      RECT 139 145 151 205 ;
      RECT 79 195 111 205 ;
      RECT 99 145 111 205 ;
      RECT 59 145 71 205 ;
      RECT 119 122.6 131 205 ;
      RECT 79 145 91 205 ;
      RECT 99 145 131 155 ;
      RECT 59 145 91 155 ;
      RECT 119 122.6 151 134.6 ;
      RECT 139 45 151 134.6 ;
    LAYER NSD ;
      RECT 260 142.25 270 190 ;
      RECT 220 142.25 230 190 ;
      RECT 180 60 190 190 ;
      RECT 180 142.25 270 152.25 ;
      RECT 90 96.35 140 106.35 ;
      RECT 130 43.35 140 106.35 ;
      RECT 90 60 100 106.35 ;
      RECT 130 43.35 183.15 53.35 ;
      RECT 130 141.75 140 190 ;
      RECT 90 141.75 100 190 ;
      RECT 50 141.75 60 190 ;
      RECT 50 141.75 140 151.75 ;
      RECT 108.6 131.2 116.6 151.75 ;
      RECT 30 96.35 80 106.35 ;
      RECT 70 42.05 80 106.35 ;
      RECT 30 60 40 106.35 ;
      RECT 110 42.05 120 90 ;
      RECT 70 42.05 120 52.05 ;
      RECT 30 160 40 190 ;
    LAYER Contact ;
      RECT 188.5 115.265 189.5 116.265 ;
      RECT 188.5 117.265 189.5 118.265 ;
      RECT 188.5 119.265 189.5 120.265 ;
      RECT 188.5 121.265 189.5 122.265 ;
      RECT 188.5 123.265 189.5 124.265 ;
      RECT 186.5 115.265 187.5 116.265 ;
      RECT 186.5 117.265 187.5 118.265 ;
      RECT 186.5 119.265 187.5 120.265 ;
      RECT 186.5 121.265 187.5 122.265 ;
      RECT 186.5 123.265 187.5 124.265 ;
      RECT 184.5 115.265 185.5 116.265 ;
      RECT 184.5 117.265 185.5 118.265 ;
      RECT 184.5 119.265 185.5 120.265 ;
      RECT 184.5 121.265 185.5 122.265 ;
      RECT 184.5 123.265 185.5 124.265 ;
      RECT 182.5 115.265 183.5 116.265 ;
      RECT 182.5 117.265 183.5 118.265 ;
      RECT 182.5 119.265 183.5 120.265 ;
      RECT 182.5 121.265 183.5 122.265 ;
      RECT 182.5 123.265 183.5 124.265 ;
      RECT 181.665 43.835 182.665 44.835 ;
      RECT 181.665 45.835 182.665 46.835 ;
      RECT 181.665 47.835 182.665 48.835 ;
      RECT 181.665 49.835 182.665 50.835 ;
      RECT 181.665 51.835 182.665 52.835 ;
      RECT 180.5 115.265 181.5 116.265 ;
      RECT 180.5 117.265 181.5 118.265 ;
      RECT 180.5 119.265 181.5 120.265 ;
      RECT 180.5 121.265 181.5 122.265 ;
      RECT 180.5 123.265 181.5 124.265 ;
      RECT 179.665 43.835 180.665 44.835 ;
      RECT 179.665 45.835 180.665 46.835 ;
      RECT 179.665 47.835 180.665 48.835 ;
      RECT 179.665 49.835 180.665 50.835 ;
      RECT 179.665 51.835 180.665 52.835 ;
      RECT 177.665 43.835 178.665 44.835 ;
      RECT 177.665 45.835 178.665 46.835 ;
      RECT 177.665 47.835 178.665 48.835 ;
      RECT 177.665 49.835 178.665 50.835 ;
      RECT 177.665 51.835 178.665 52.835 ;
      RECT 175.665 43.835 176.665 44.835 ;
      RECT 175.665 45.835 176.665 46.835 ;
      RECT 175.665 47.835 176.665 48.835 ;
      RECT 175.665 49.835 176.665 50.835 ;
      RECT 175.665 51.835 176.665 52.835 ;
      RECT 173.665 43.835 174.665 44.835 ;
      RECT 173.665 45.835 174.665 46.835 ;
      RECT 173.665 47.835 174.665 48.835 ;
      RECT 173.665 49.835 174.665 50.835 ;
      RECT 173.665 51.835 174.665 52.835 ;
      RECT 115.11 131.675 116.11 132.675 ;
      RECT 115.11 133.675 116.11 134.675 ;
      RECT 115.11 135.675 116.11 136.675 ;
      RECT 115.11 137.675 116.11 138.675 ;
      RECT 113.11 131.675 114.11 132.675 ;
      RECT 113.11 133.675 114.11 134.675 ;
      RECT 113.11 135.675 114.11 136.675 ;
      RECT 113.11 137.675 114.11 138.675 ;
      RECT 111.11 131.675 112.11 132.675 ;
      RECT 111.11 133.675 112.11 134.675 ;
      RECT 111.11 135.675 112.11 136.675 ;
      RECT 111.11 137.675 112.11 138.675 ;
      RECT 109.11 131.675 110.11 132.675 ;
      RECT 109.11 133.675 110.11 134.675 ;
      RECT 109.11 135.675 110.11 136.675 ;
      RECT 109.11 137.675 110.11 138.675 ;
    LAYER Cont ;
      RECT 203.5 115.265 204.5 116.265 ;
      RECT 203.5 117.265 204.5 118.265 ;
      RECT 203.5 119.265 204.5 120.265 ;
      RECT 203.5 121.265 204.5 122.265 ;
      RECT 203.5 123.265 204.5 124.265 ;
      RECT 201.5 115.265 202.5 116.265 ;
      RECT 201.5 117.265 202.5 118.265 ;
      RECT 201.5 119.265 202.5 120.265 ;
      RECT 201.5 121.265 202.5 122.265 ;
      RECT 201.5 123.265 202.5 124.265 ;
      RECT 199.5 115.265 200.5 116.265 ;
      RECT 199.5 117.265 200.5 118.265 ;
      RECT 199.5 119.265 200.5 120.265 ;
      RECT 199.5 121.265 200.5 122.265 ;
      RECT 199.5 123.265 200.5 124.265 ;
      RECT 197.5 43.835 198.5 44.835 ;
      RECT 197.5 45.835 198.5 46.835 ;
      RECT 197.5 47.835 198.5 48.835 ;
      RECT 197.5 49.835 198.5 50.835 ;
      RECT 197.5 51.835 198.5 52.835 ;
      RECT 197.5 115.265 198.5 116.265 ;
      RECT 197.5 117.265 198.5 118.265 ;
      RECT 197.5 119.265 198.5 120.265 ;
      RECT 197.5 121.265 198.5 122.265 ;
      RECT 197.5 123.265 198.5 124.265 ;
      RECT 195.5 43.835 196.5 44.835 ;
      RECT 195.5 45.835 196.5 46.835 ;
      RECT 195.5 47.835 196.5 48.835 ;
      RECT 195.5 49.835 196.5 50.835 ;
      RECT 195.5 51.835 196.5 52.835 ;
      RECT 195.5 115.265 196.5 116.265 ;
      RECT 195.5 117.265 196.5 118.265 ;
      RECT 195.5 119.265 196.5 120.265 ;
      RECT 195.5 121.265 196.5 122.265 ;
      RECT 195.5 123.265 196.5 124.265 ;
      RECT 193.5 43.835 194.5 44.835 ;
      RECT 193.5 45.835 194.5 46.835 ;
      RECT 193.5 47.835 194.5 48.835 ;
      RECT 193.5 49.835 194.5 50.835 ;
      RECT 193.5 51.835 194.5 52.835 ;
      RECT 191.5 43.835 192.5 44.835 ;
      RECT 191.5 45.835 192.5 46.835 ;
      RECT 191.5 47.835 192.5 48.835 ;
      RECT 191.5 49.835 192.5 50.835 ;
      RECT 191.5 51.835 192.5 52.835 ;
      RECT 189.5 43.835 190.5 44.835 ;
      RECT 189.5 45.835 190.5 46.835 ;
      RECT 189.5 47.835 190.5 48.835 ;
      RECT 189.5 49.835 190.5 50.835 ;
      RECT 189.5 51.835 190.5 52.835 ;
      RECT 126.925 131.675 127.925 132.675 ;
      RECT 126.925 133.675 127.925 134.675 ;
      RECT 126.925 135.675 127.925 136.675 ;
      RECT 126.925 137.675 127.925 138.675 ;
      RECT 124.925 131.675 125.925 132.675 ;
      RECT 124.925 133.675 125.925 134.675 ;
      RECT 124.925 135.675 125.925 136.675 ;
      RECT 124.925 137.675 125.925 138.675 ;
      RECT 122.925 131.675 123.925 132.675 ;
      RECT 122.925 133.675 123.925 134.675 ;
      RECT 122.925 135.675 123.925 136.675 ;
      RECT 122.925 137.675 123.925 138.675 ;
      RECT 120.925 131.675 121.925 132.675 ;
      RECT 120.925 133.675 121.925 134.675 ;
      RECT 120.925 135.675 121.925 136.675 ;
      RECT 120.925 137.675 121.925 138.675 ;
    LAYER Metal1 ;
      RECT 180 114.765 205 124.765 ;
      RECT 173.165 43.335 199 53.335 ;
      RECT 108.61 131.175 128.425 139.175 ;
  END
END MoS2And

MACRO MoS2DFlipFlop
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MoS2DFlipFlop 0 0 ;
  SIZE 1300 BY 280 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN CP
    DIRECTION INOUT ;
    USE CLOCK ;
    PORT
      LAYER Gate ;
        RECT 799 25.9 811 135.05 ;
        RECT 539 25.9 811 33.9 ;
        RECT 719 25.9 731 135.05 ;
        RECT 539 25.9 551 105 ;
        RECT 519 45 551 55 ;
        RECT 479 122 531 134 ;
        RECT 519 45 531 134 ;
        RECT 479 122 491 205 ;
      LAYER Metal1 ;
        RECT 469.452 196.748 488.152 204.748 ;
      LAYER NSD ;
        RECT 469.452 196.748 477.452 204.748 ;
      LAYER Cont ;
        RECT 480.652 203.248 481.652 204.248 ;
        RECT 480.652 201.248 481.652 202.248 ;
        RECT 480.652 199.248 481.652 200.248 ;
        RECT 480.652 197.248 481.652 198.248 ;
        RECT 482.652 203.248 483.652 204.248 ;
        RECT 482.652 201.248 483.652 202.248 ;
        RECT 482.652 199.248 483.652 200.248 ;
        RECT 482.652 197.248 483.652 198.248 ;
        RECT 484.652 203.248 485.652 204.248 ;
        RECT 484.652 201.248 485.652 202.248 ;
        RECT 484.652 199.248 485.652 200.248 ;
        RECT 484.652 197.248 485.652 198.248 ;
        RECT 486.652 203.248 487.652 204.248 ;
        RECT 486.652 201.248 487.652 202.248 ;
        RECT 486.652 199.248 487.652 200.248 ;
        RECT 486.652 197.248 487.652 198.248 ;
      LAYER Contact ;
        RECT 469.952 203.248 470.952 204.248 ;
        RECT 469.952 201.248 470.952 202.248 ;
        RECT 469.952 199.248 470.952 200.248 ;
        RECT 469.952 197.248 470.952 198.248 ;
        RECT 471.952 203.248 472.952 204.248 ;
        RECT 471.952 201.248 472.952 202.248 ;
        RECT 471.952 199.248 472.952 200.248 ;
        RECT 471.952 197.248 472.952 198.248 ;
        RECT 473.952 203.248 474.952 204.248 ;
        RECT 473.952 201.248 474.952 202.248 ;
        RECT 473.952 199.248 474.952 200.248 ;
        RECT 473.952 197.248 474.952 198.248 ;
        RECT 475.952 203.248 476.952 204.248 ;
        RECT 475.952 201.248 476.952 202.248 ;
        RECT 475.952 199.248 476.952 200.248 ;
        RECT 475.952 197.248 476.952 198.248 ;
    END
  END CP
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 99 45 111 105 ;
        RECT 79 45 111 55 ;
        RECT 39 122 91 134 ;
        RECT 79 45 91 134 ;
        RECT 39 122 51 205 ;
      LAYER Metal1 ;
        RECT 40.696 196.628 48.696 215.852 ;
      LAYER NSD ;
        RECT 40.696 207.852 48.696 215.852 ;
      LAYER Cont ;
        RECT 41.196 203.128 42.196 204.128 ;
        RECT 41.196 201.128 42.196 202.128 ;
        RECT 41.196 199.128 42.196 200.128 ;
        RECT 41.196 197.128 42.196 198.128 ;
        RECT 43.196 203.128 44.196 204.128 ;
        RECT 43.196 201.128 44.196 202.128 ;
        RECT 43.196 199.128 44.196 200.128 ;
        RECT 43.196 197.128 44.196 198.128 ;
        RECT 45.196 203.128 46.196 204.128 ;
        RECT 45.196 201.128 46.196 202.128 ;
        RECT 45.196 199.128 46.196 200.128 ;
        RECT 45.196 197.128 46.196 198.128 ;
        RECT 47.196 203.128 48.196 204.128 ;
        RECT 47.196 201.128 48.196 202.128 ;
        RECT 47.196 199.128 48.196 200.128 ;
        RECT 47.196 197.128 48.196 198.128 ;
      LAYER Contact ;
        RECT 41.196 214.352 42.196 215.352 ;
        RECT 41.196 212.352 42.196 213.352 ;
        RECT 41.196 210.352 42.196 211.352 ;
        RECT 41.196 208.352 42.196 209.352 ;
        RECT 43.196 214.352 44.196 215.352 ;
        RECT 43.196 212.352 44.196 213.352 ;
        RECT 43.196 210.352 44.196 211.352 ;
        RECT 43.196 208.352 44.196 209.352 ;
        RECT 45.196 214.352 46.196 215.352 ;
        RECT 45.196 212.352 46.196 213.352 ;
        RECT 45.196 210.352 46.196 211.352 ;
        RECT 45.196 208.352 46.196 209.352 ;
        RECT 47.196 214.352 48.196 215.352 ;
        RECT 47.196 212.352 48.196 213.352 ;
        RECT 47.196 210.352 48.196 211.352 ;
        RECT 47.196 208.352 48.196 209.352 ;
    END
  END D
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 10 0 20 190 ;
    END
    PORT
      LAYER NSD ;
        RECT 50 0 60 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 230 0 240 190 ;
    END
    PORT
      LAYER NSD ;
        RECT 270 0 280 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 450 0 460 190 ;
    END
    PORT
      LAYER NSD ;
        RECT 490 0 500 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 670 0 680 134.05 ;
    END
    PORT
      LAYER NSD ;
        RECT 750 0 760 134.05 ;
    END
    PORT
      LAYER NSD ;
        RECT 870 0 880 190 ;
    END
    PORT
      LAYER NSD ;
        RECT 870 44.35 920 54.35 ;
    END
    PORT
      LAYER NSD ;
        RECT 910 44.35 920 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 1090 0 1100 190 ;
    END
    PORT
      LAYER NSD ;
        RECT 1090 43.45 1140 53.45 ;
    END
    PORT
      LAYER NSD ;
        RECT 1130 43.45 1140 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 0 1300 20 ;
    END
  END GND
  PIN NQ
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 899 32.7 1208.95 40.7 ;
        RECT 899 32.7 911 105 ;
        RECT 879 45 911 55 ;
        RECT 879 45 891 205 ;
      LAYER Metal1 ;
        RECT 1200.58 32.68 1218.696 40.68 ;
      LAYER NSD ;
        RECT 1170 96.35 1220 106.35 ;
        RECT 1210 31.7 1220 106.35 ;
        RECT 1170 60 1180 106.35 ;
      LAYER Cont ;
        RECT 1201.08 39.18 1202.08 40.18 ;
        RECT 1201.08 37.18 1202.08 38.18 ;
        RECT 1201.08 35.18 1202.08 36.18 ;
        RECT 1201.08 33.18 1202.08 34.18 ;
        RECT 1203.08 39.18 1204.08 40.18 ;
        RECT 1203.08 37.18 1204.08 38.18 ;
        RECT 1203.08 35.18 1204.08 36.18 ;
        RECT 1203.08 33.18 1204.08 34.18 ;
        RECT 1205.08 39.18 1206.08 40.18 ;
        RECT 1205.08 37.18 1206.08 38.18 ;
        RECT 1205.08 35.18 1206.08 36.18 ;
        RECT 1205.08 33.18 1206.08 34.18 ;
        RECT 1207.08 39.18 1208.08 40.18 ;
        RECT 1207.08 37.18 1208.08 38.18 ;
        RECT 1207.08 35.18 1208.08 36.18 ;
        RECT 1207.08 33.18 1208.08 34.18 ;
      LAYER Contact ;
        RECT 1211.196 39.18 1212.196 40.18 ;
        RECT 1211.196 37.18 1212.196 38.18 ;
        RECT 1211.196 35.18 1212.196 36.18 ;
        RECT 1211.196 33.18 1212.196 34.18 ;
        RECT 1213.196 39.18 1214.196 40.18 ;
        RECT 1213.196 37.18 1214.196 38.18 ;
        RECT 1213.196 35.18 1214.196 36.18 ;
        RECT 1213.196 33.18 1214.196 34.18 ;
        RECT 1215.196 39.18 1216.196 40.18 ;
        RECT 1215.196 37.18 1216.196 38.18 ;
        RECT 1215.196 35.18 1216.196 36.18 ;
        RECT 1215.196 33.18 1216.196 34.18 ;
        RECT 1217.196 39.18 1218.196 40.18 ;
        RECT 1217.196 37.18 1218.196 38.18 ;
        RECT 1217.196 35.18 1218.196 36.18 ;
        RECT 1217.196 33.18 1218.196 34.18 ;
    END
  END NQ
  PIN Q
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 1179 45 1191 105 ;
        RECT 1159 45 1191 55 ;
        RECT 1119 122 1171 134 ;
        RECT 1159 45 1171 134 ;
        RECT 1119 122 1131 205 ;
      LAYER Metal1 ;
        RECT 1077.4 124.25 1127.35 132.25 ;
        RECT 1077.4 97.05 1085.4 132.25 ;
        RECT 989.4 97.05 1085.4 105.05 ;
      LAYER NSD ;
        RECT 950 96.35 1000 106.35 ;
        RECT 990 60 1000 106.35 ;
        RECT 950 60 960 106.35 ;
      LAYER Cont ;
        RECT 1119.872 130.772 1120.872 131.772 ;
        RECT 1119.872 128.772 1120.872 129.772 ;
        RECT 1119.872 126.772 1120.872 127.772 ;
        RECT 1119.872 124.772 1120.872 125.772 ;
        RECT 1121.872 130.772 1122.872 131.772 ;
        RECT 1121.872 128.772 1122.872 129.772 ;
        RECT 1121.872 126.772 1122.872 127.772 ;
        RECT 1121.872 124.772 1122.872 125.772 ;
        RECT 1123.872 130.772 1124.872 131.772 ;
        RECT 1123.872 128.772 1124.872 129.772 ;
        RECT 1123.872 126.772 1124.872 127.772 ;
        RECT 1123.872 124.772 1124.872 125.772 ;
        RECT 1125.872 130.772 1126.872 131.772 ;
        RECT 1125.872 128.772 1126.872 129.772 ;
        RECT 1125.872 126.772 1126.872 127.772 ;
        RECT 1125.872 124.772 1126.872 125.772 ;
      LAYER Contact ;
        RECT 989.916 103.532 990.916 104.532 ;
        RECT 989.916 101.532 990.916 102.532 ;
        RECT 989.916 99.532 990.916 100.532 ;
        RECT 989.916 97.532 990.916 98.532 ;
        RECT 991.916 103.532 992.916 104.532 ;
        RECT 991.916 101.532 992.916 102.532 ;
        RECT 991.916 99.532 992.916 100.532 ;
        RECT 991.916 97.532 992.916 98.532 ;
        RECT 993.916 103.532 994.916 104.532 ;
        RECT 993.916 101.532 994.916 102.532 ;
        RECT 993.916 99.532 994.916 100.532 ;
        RECT 993.916 97.532 994.916 98.532 ;
        RECT 995.916 103.532 996.916 104.532 ;
        RECT 995.916 101.532 996.916 102.532 ;
        RECT 995.916 99.532 996.916 100.532 ;
        RECT 995.916 97.532 996.916 98.532 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Contact ;
        RECT 1255.4 212.916 1256.4 213.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1255.4 214.916 1256.4 215.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1255.4 216.916 1256.4 217.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1255.4 218.916 1256.4 219.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1255.4 261.912 1256.4 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1255.4 263.912 1256.4 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1255.4 265.912 1256.4 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1255.4 267.912 1256.4 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1253.4 212.916 1254.4 213.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1253.4 214.916 1254.4 215.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1253.4 216.916 1254.4 217.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1253.4 218.916 1254.4 219.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1253.4 261.912 1254.4 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1253.4 263.912 1254.4 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1253.4 265.912 1254.4 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1253.4 267.912 1254.4 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1251.4 212.916 1252.4 213.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1251.4 214.916 1252.4 215.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1251.4 216.916 1252.4 217.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1251.4 218.916 1252.4 219.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1251.4 261.912 1252.4 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1251.4 263.912 1252.4 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1251.4 265.912 1252.4 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1251.4 267.912 1252.4 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1249.4 212.916 1250.4 213.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1249.4 214.916 1250.4 215.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1249.4 216.916 1250.4 217.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1249.4 218.916 1250.4 219.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1249.4 261.912 1250.4 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1249.4 263.912 1250.4 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1249.4 265.912 1250.4 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1249.4 267.912 1250.4 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1035.868 212.916 1036.868 213.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1035.868 214.916 1036.868 215.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1035.868 216.916 1036.868 217.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1035.868 218.916 1036.868 219.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1035.868 261.912 1036.868 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1035.868 263.912 1036.868 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1035.868 265.912 1036.868 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1035.868 267.912 1036.868 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1033.868 212.916 1034.868 213.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1033.868 214.916 1034.868 215.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1033.868 216.916 1034.868 217.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1033.868 218.916 1034.868 219.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1033.868 261.912 1034.868 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1033.868 263.912 1034.868 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1033.868 265.912 1034.868 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1033.868 267.912 1034.868 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1031.868 212.916 1032.868 213.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1031.868 214.916 1032.868 215.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1031.868 216.916 1032.868 217.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1031.868 218.916 1032.868 219.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1031.868 261.912 1032.868 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1031.868 263.912 1032.868 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1031.868 265.912 1032.868 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1031.868 267.912 1032.868 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1029.868 212.916 1030.868 213.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1029.868 214.916 1030.868 215.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1029.868 216.916 1030.868 217.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1029.868 218.916 1030.868 219.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 1029.868 261.912 1030.868 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1029.868 263.912 1030.868 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1029.868 265.912 1030.868 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 1029.868 267.912 1030.868 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 797.336 216.06 798.336 217.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 797.336 218.06 798.336 219.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 797.336 220.06 798.336 221.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 797.336 222.06 798.336 223.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 797.336 262.116 798.336 263.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 797.336 264.116 798.336 265.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 797.336 266.116 798.336 267.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 797.336 268.116 798.336 269.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 795.336 216.06 796.336 217.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 795.336 218.06 796.336 219.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 795.336 220.06 796.336 221.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 795.336 222.06 796.336 223.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 795.336 262.116 796.336 263.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 795.336 264.116 796.336 265.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 795.336 266.116 796.336 267.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 795.336 268.116 796.336 269.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 793.336 216.06 794.336 217.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 793.336 218.06 794.336 219.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 793.336 220.06 794.336 221.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 793.336 222.06 794.336 223.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 793.336 262.116 794.336 263.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 793.336 264.116 794.336 265.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 793.336 266.116 794.336 267.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 793.336 268.116 794.336 269.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 791.336 216.06 792.336 217.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 791.336 218.06 792.336 219.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 791.336 220.06 792.336 221.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 791.336 222.06 792.336 223.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 791.336 262.116 792.336 263.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 791.336 264.116 792.336 265.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 791.336 266.116 792.336 267.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 791.336 268.116 792.336 269.116 ;
    END
    PORT
      LAYER Contact ;
        RECT 613.568 219.536 614.568 220.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 613.568 221.536 614.568 222.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 613.568 223.536 614.568 224.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 613.568 225.536 614.568 226.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 613.568 261.912 614.568 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 613.568 263.912 614.568 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 613.568 265.912 614.568 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 613.568 267.912 614.568 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 611.568 219.536 612.568 220.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 611.568 221.536 612.568 222.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 611.568 223.536 612.568 224.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 611.568 225.536 612.568 226.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 611.568 261.912 612.568 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 611.568 263.912 612.568 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 611.568 265.912 612.568 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 611.568 267.912 612.568 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 609.568 219.536 610.568 220.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 609.568 221.536 610.568 222.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 609.568 223.536 610.568 224.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 609.568 225.536 610.568 226.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 609.568 261.912 610.568 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 609.568 263.912 610.568 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 609.568 265.912 610.568 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 609.568 267.912 610.568 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 607.568 219.536 608.568 220.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 607.568 221.536 608.568 222.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 607.568 223.536 608.568 224.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 607.568 225.536 608.568 226.536 ;
    END
    PORT
      LAYER Contact ;
        RECT 607.568 261.912 608.568 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 607.568 263.912 608.568 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 607.568 265.912 608.568 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 607.568 267.912 608.568 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 395.296 219.356 396.296 220.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 395.296 221.356 396.296 222.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 395.296 223.356 396.296 224.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 395.296 225.356 396.296 226.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 395.296 261.912 396.296 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 395.296 263.912 396.296 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 395.296 265.912 396.296 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 395.296 267.912 396.296 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 393.296 219.356 394.296 220.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 393.296 221.356 394.296 222.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 393.296 223.356 394.296 224.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 393.296 225.356 394.296 226.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 393.296 261.912 394.296 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 393.296 263.912 394.296 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 393.296 265.912 394.296 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 393.296 267.912 394.296 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 391.296 219.356 392.296 220.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 391.296 221.356 392.296 222.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 391.296 223.356 392.296 224.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 391.296 225.356 392.296 226.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 391.296 261.912 392.296 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 391.296 263.912 392.296 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 391.296 265.912 392.296 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 391.296 267.912 392.296 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 389.296 219.356 390.296 220.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 389.296 221.356 390.296 222.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 389.296 223.356 390.296 224.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 389.296 225.356 390.296 226.356 ;
    END
    PORT
      LAYER Contact ;
        RECT 389.296 261.912 390.296 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 389.296 263.912 390.296 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 389.296 265.912 390.296 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 389.296 267.912 390.296 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 175.656 212.916 176.656 213.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 175.656 214.916 176.656 215.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 175.656 216.916 176.656 217.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 175.656 218.916 176.656 219.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 175.656 261.912 176.656 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 175.656 263.912 176.656 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 175.656 265.912 176.656 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 175.656 267.912 176.656 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.656 212.916 174.656 213.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.656 214.916 174.656 215.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.656 216.916 174.656 217.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.656 218.916 174.656 219.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.656 261.912 174.656 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.656 263.912 174.656 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.656 265.912 174.656 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.656 267.912 174.656 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.656 212.916 172.656 213.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.656 214.916 172.656 215.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.656 216.916 172.656 217.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.656 218.916 172.656 219.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.656 261.912 172.656 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.656 263.912 172.656 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.656 265.912 172.656 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.656 267.912 172.656 268.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.656 212.916 170.656 213.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.656 214.916 170.656 215.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.656 216.916 170.656 217.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.656 218.916 170.656 219.916 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.656 261.912 170.656 262.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.656 263.912 170.656 264.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.656 265.912 170.656 266.912 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.656 267.912 170.656 268.912 ;
    END
    PORT
      LAYER NSD ;
        RECT 150 60 160 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 150 98.9 178.25 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 168.25 98.9 178.25 220.75 ;
    END
    PORT
      LAYER NSD ;
        RECT 370 60 380 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 370 98.9 397.95 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 387.95 98.9 397.95 226.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 590 60 600 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 590 98.9 616.2 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 606.2 98.9 616.2 227.05 ;
    END
    PORT
      LAYER NSD ;
        RECT 790 170 800 223.58 ;
    END
    PORT
      LAYER NSD ;
        RECT 1010 60 1020 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 1010 98.9 1038.35 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 1028.35 98.9 1038.35 220.75 ;
    END
    PORT
      LAYER NSD ;
        RECT 1230 60 1240 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 1230 98.9 1257.65 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 1247.65 98.9 1257.65 220.75 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 260 1300 280 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 169.156 212.416 177.156 269.412 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 388.796 218.856 396.796 269.412 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 607.068 219.036 615.068 269.412 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 790.836 215.56 798.836 269.616 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 1029.368 212.416 1037.368 269.412 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 1248.9 212.416 1256.9 269.412 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 70 160 80 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 110 160 120 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 150 160 160 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 70 198.1 160 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 290 160 300 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 330 160 340 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 370 160 380 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 290 198.1 380 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 510 160 520 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 550 160 560 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 590 160 600 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 510 198.1 600 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 690 170 700 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 730 170 740 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 770 170 780 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 930 160 940 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 970 160 980 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 1010 160 1020 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 930 198.1 1020 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 1150 160 1160 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 1190 160 1200 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 1230 160 1240 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 1150 198.1 1240 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 230 1300 250 ;
    END
  END VSS
  OBS
    LAYER Gate ;
      RECT 1199 195 1231 205 ;
      RECT 1219 145 1231 205 ;
      RECT 1159 195 1191 205 ;
      RECT 1179 145 1191 205 ;
      RECT 1139 145 1151 205 ;
      RECT 1199 122.6 1211 205 ;
      RECT 1159 145 1171 205 ;
      RECT 1179 145 1211 155 ;
      RECT 1139 145 1171 155 ;
      RECT 1199 122.6 1231 134.6 ;
      RECT 1219 45 1231 134.6 ;
      RECT 1099 45 1111 205 ;
      RECT 1119 45 1131 105 ;
      RECT 1099 45 1131 55 ;
      RECT 979 195 1011 205 ;
      RECT 999 145 1011 205 ;
      RECT 939 195 971 205 ;
      RECT 959 145 971 205 ;
      RECT 919 145 931 205 ;
      RECT 979 122.6 991 205 ;
      RECT 939 145 951 205 ;
      RECT 959 145 991 155 ;
      RECT 919 145 951 155 ;
      RECT 979 122.6 1011 134.6 ;
      RECT 999 45 1011 134.6 ;
      RECT 899 122 911 195 ;
      RECT 899 122 951 134 ;
      RECT 939 45 951 134 ;
      RECT 959 45 971 105 ;
      RECT 939 45 971 55 ;
      RECT 739 205 771 215 ;
      RECT 759 155 771 215 ;
      RECT 699 205 731 215 ;
      RECT 719 155 731 215 ;
      RECT 679 155 691 215 ;
      RECT 799 155 811 205.1 ;
      RECT 739 155 751 215 ;
      RECT 699 155 711 215 ;
      RECT 759 155 811 167 ;
      RECT 719 155 751 165 ;
      RECT 679 155 711 165 ;
      RECT 779 43.05 791 135.05 ;
      RECT 781.15 35.2 789.15 135.05 ;
      RECT 679 138 771 146 ;
      RECT 759 43.25 771 146 ;
      RECT 679 43.45 691 146 ;
      RECT 699 43.05 711 135.05 ;
      RECT 701.25 35.2 709.25 135.05 ;
      RECT 259 209.6 650.35 217.6 ;
      RECT 259 122 271 217.6 ;
      RECT 259 122 311 134 ;
      RECT 299 45 311 134 ;
      RECT 319 45 331 105 ;
      RECT 299 45 331 55 ;
      RECT 559 195 591 205 ;
      RECT 579 145 591 205 ;
      RECT 519 195 551 205 ;
      RECT 539 145 551 205 ;
      RECT 499 145 511 205 ;
      RECT 559 122.6 571 205 ;
      RECT 519 145 531 205 ;
      RECT 539 145 571 155 ;
      RECT 499 145 531 155 ;
      RECT 559 122.6 591 134.6 ;
      RECT 579 45 591 134.6 ;
      RECT 19 45 31 205 ;
      RECT 39 33.75 51 105 ;
      RECT 19 45 51 55 ;
      RECT 39 33.75 529.8 41.75 ;
      RECT 521.8 25.05 529.8 41.75 ;
      RECT 459 45 471 195 ;
      RECT 479 45 491 105 ;
      RECT 459 45 491 55 ;
      RECT 363.85 45 491 53 ;
      RECT 339 195 371 205 ;
      RECT 359 145 371 205 ;
      RECT 299 195 331 205 ;
      RECT 319 145 331 205 ;
      RECT 279 145 291 205 ;
      RECT 339 122.6 351 205 ;
      RECT 299 145 311 205 ;
      RECT 319 145 351 155 ;
      RECT 279 145 311 155 ;
      RECT 339 122.6 371 134.6 ;
      RECT 359 55 371 134.6 ;
      RECT 239 45 251 205 ;
      RECT 259 45 271 105 ;
      RECT 239 45 271 55 ;
      RECT 142.85 45 271 53 ;
      RECT 119 195 151 205 ;
      RECT 139 145 151 205 ;
      RECT 79 195 111 205 ;
      RECT 99 145 111 205 ;
      RECT 59 145 71 205 ;
      RECT 119 122.6 131 205 ;
      RECT 79 145 91 205 ;
      RECT 99 145 131 155 ;
      RECT 59 145 91 155 ;
      RECT 119 122.6 151 134.6 ;
      RECT 139 55 151 134.6 ;
    LAYER NSD ;
      RECT 1210 141.75 1220 190 ;
      RECT 1170 141.75 1180 190 ;
      RECT 1130 141.75 1140 190 ;
      RECT 1130 141.75 1220 151.75 ;
      RECT 1188.6 131.2 1196.6 151.75 ;
      RECT 1110 96.35 1160 106.35 ;
      RECT 1150 44.85 1160 106.35 ;
      RECT 1110 60 1120 106.35 ;
      RECT 1190 44.85 1200 90 ;
      RECT 1150 44.85 1200 54.85 ;
      RECT 990 141.75 1000 190 ;
      RECT 950 141.75 960 190 ;
      RECT 910 141.75 920 190 ;
      RECT 910 141.75 1000 151.75 ;
      RECT 968.6 131.2 976.6 151.75 ;
      RECT 890 96.35 940 106.35 ;
      RECT 930 45.1 940 106.35 ;
      RECT 890 60 900 106.35 ;
      RECT 970 45.1 980 90 ;
      RECT 930 45.1 980 55.1 ;
      RECT 810 27.75 820 200 ;
      RECT 812 25.05 820 200 ;
      RECT 670 154.5 680 215.25 ;
      RECT 750 154.5 760 200 ;
      RECT 710 154.5 720 200 ;
      RECT 670 154.5 760 164.5 ;
      RECT 730 44.05 740 164.5 ;
      RECT 530 96.35 580 106.35 ;
      RECT 570 60 580 106.35 ;
      RECT 530 60 540 106.35 ;
      RECT 570 141.75 580 190 ;
      RECT 530 141.75 540 190 ;
      RECT 490 141.75 500 190 ;
      RECT 490 141.75 580 151.75 ;
      RECT 548.6 131.2 556.6 151.75 ;
      RECT 470 96.35 520 106.35 ;
      RECT 510 46.8 520 106.35 ;
      RECT 470 60 480 106.35 ;
      RECT 550 46.8 560 90 ;
      RECT 510 46.8 560 56.8 ;
      RECT 310 96.35 360 106.35 ;
      RECT 350 44 360 106.35 ;
      RECT 310 60 320 106.35 ;
      RECT 350 141.75 360 190 ;
      RECT 310 141.75 320 190 ;
      RECT 270 141.75 280 190 ;
      RECT 270 141.75 360 151.75 ;
      RECT 328.6 131.2 336.6 151.75 ;
      RECT 250 96.35 300 106.35 ;
      RECT 290 42.05 300 106.35 ;
      RECT 250 60 260 106.35 ;
      RECT 330 42.05 340 90 ;
      RECT 290 42.05 340 52.05 ;
      RECT 90 96.35 140 106.35 ;
      RECT 130 44 140 106.35 ;
      RECT 90 60 100 106.35 ;
      RECT 130 141.75 140 190 ;
      RECT 90 141.75 100 190 ;
      RECT 50 141.75 60 190 ;
      RECT 50 141.75 140 151.75 ;
      RECT 108.6 131.2 116.6 151.75 ;
      RECT 30 96.35 80 106.35 ;
      RECT 70 42.05 80 106.35 ;
      RECT 30 60 40 106.35 ;
      RECT 110 42.05 120 90 ;
      RECT 70 42.05 120 52.05 ;
      RECT 1110 160 1120 190 ;
      RECT 890 160 900 190 ;
      RECT 790 44.032 800 134.032 ;
      RECT 770 44.032 780 134.032 ;
      RECT 710 44.032 720 134.032 ;
      RECT 690 44.032 700 134.032 ;
      RECT 651.388 97.176 659.388 217.596 ;
      RECT 470 160 480 190 ;
      RECT 250 160 260 190 ;
      RECT 30 160 40 190 ;
    LAYER Contact ;
      RECT 1195.112 131.676 1196.112 132.676 ;
      RECT 1195.112 133.676 1196.112 134.676 ;
      RECT 1195.112 135.676 1196.112 136.676 ;
      RECT 1195.112 137.676 1196.112 138.676 ;
      RECT 1193.112 131.676 1194.112 132.676 ;
      RECT 1193.112 133.676 1194.112 134.676 ;
      RECT 1193.112 135.676 1194.112 136.676 ;
      RECT 1193.112 137.676 1194.112 138.676 ;
      RECT 1191.112 131.676 1192.112 132.676 ;
      RECT 1191.112 133.676 1192.112 134.676 ;
      RECT 1191.112 135.676 1192.112 136.676 ;
      RECT 1191.112 137.676 1192.112 138.676 ;
      RECT 1189.112 131.676 1190.112 132.676 ;
      RECT 1189.112 133.676 1190.112 134.676 ;
      RECT 1189.112 135.676 1190.112 136.676 ;
      RECT 1189.112 137.676 1190.112 138.676 ;
      RECT 975.112 131.676 976.112 132.676 ;
      RECT 975.112 133.676 976.112 134.676 ;
      RECT 975.112 135.676 976.112 136.676 ;
      RECT 975.112 137.676 976.112 138.676 ;
      RECT 973.112 131.676 974.112 132.676 ;
      RECT 973.112 133.676 974.112 134.676 ;
      RECT 973.112 135.676 974.112 136.676 ;
      RECT 973.112 137.676 974.112 138.676 ;
      RECT 971.112 131.676 972.112 132.676 ;
      RECT 971.112 133.676 972.112 134.676 ;
      RECT 971.112 135.676 972.112 136.676 ;
      RECT 971.112 137.676 972.112 138.676 ;
      RECT 969.112 131.676 970.112 132.676 ;
      RECT 969.112 133.676 970.112 134.676 ;
      RECT 969.112 135.676 970.112 136.676 ;
      RECT 969.112 137.676 970.112 138.676 ;
      RECT 818.5 25.536 819.5 26.536 ;
      RECT 818.5 27.536 819.5 28.536 ;
      RECT 818.5 29.536 819.5 30.536 ;
      RECT 818.5 31.536 819.5 32.536 ;
      RECT 816.5 25.536 817.5 26.536 ;
      RECT 816.5 27.536 817.5 28.536 ;
      RECT 816.5 29.536 817.5 30.536 ;
      RECT 816.5 31.536 817.5 32.536 ;
      RECT 814.5 25.536 815.5 26.536 ;
      RECT 814.5 27.536 815.5 28.536 ;
      RECT 814.5 29.536 815.5 30.536 ;
      RECT 814.5 31.536 815.5 32.536 ;
      RECT 812.5 25.536 813.5 26.536 ;
      RECT 812.5 27.536 813.5 28.536 ;
      RECT 812.5 29.536 813.5 30.536 ;
      RECT 812.5 31.536 813.5 32.536 ;
      RECT 676.556 206.772 677.556 207.772 ;
      RECT 676.556 208.772 677.556 209.772 ;
      RECT 676.556 210.772 677.556 211.772 ;
      RECT 676.556 212.772 677.556 213.772 ;
      RECT 674.556 206.772 675.556 207.772 ;
      RECT 674.556 208.772 675.556 209.772 ;
      RECT 674.556 210.772 675.556 211.772 ;
      RECT 674.556 212.772 675.556 213.772 ;
      RECT 672.556 206.772 673.556 207.772 ;
      RECT 672.556 208.772 673.556 209.772 ;
      RECT 672.556 210.772 673.556 211.772 ;
      RECT 672.556 212.772 673.556 213.772 ;
      RECT 670.556 206.772 671.556 207.772 ;
      RECT 670.556 208.772 671.556 209.772 ;
      RECT 670.556 210.772 671.556 211.772 ;
      RECT 670.556 212.772 671.556 213.772 ;
      RECT 657.888 97.676 658.888 98.676 ;
      RECT 657.888 99.676 658.888 100.676 ;
      RECT 657.888 101.676 658.888 102.676 ;
      RECT 657.888 103.676 658.888 104.676 ;
      RECT 657.888 138.5 658.888 139.5 ;
      RECT 657.888 140.5 658.888 141.5 ;
      RECT 657.888 142.5 658.888 143.5 ;
      RECT 657.888 144.5 658.888 145.5 ;
      RECT 657.888 210.096 658.888 211.096 ;
      RECT 657.888 212.096 658.888 213.096 ;
      RECT 657.888 214.096 658.888 215.096 ;
      RECT 657.888 216.096 658.888 217.096 ;
      RECT 655.888 97.676 656.888 98.676 ;
      RECT 655.888 99.676 656.888 100.676 ;
      RECT 655.888 101.676 656.888 102.676 ;
      RECT 655.888 103.676 656.888 104.676 ;
      RECT 655.888 138.5 656.888 139.5 ;
      RECT 655.888 140.5 656.888 141.5 ;
      RECT 655.888 142.5 656.888 143.5 ;
      RECT 655.888 144.5 656.888 145.5 ;
      RECT 655.888 210.096 656.888 211.096 ;
      RECT 655.888 212.096 656.888 213.096 ;
      RECT 655.888 214.096 656.888 215.096 ;
      RECT 655.888 216.096 656.888 217.096 ;
      RECT 653.888 97.676 654.888 98.676 ;
      RECT 653.888 99.676 654.888 100.676 ;
      RECT 653.888 101.676 654.888 102.676 ;
      RECT 653.888 103.676 654.888 104.676 ;
      RECT 653.888 138.5 654.888 139.5 ;
      RECT 653.888 140.5 654.888 141.5 ;
      RECT 653.888 142.5 654.888 143.5 ;
      RECT 653.888 144.5 654.888 145.5 ;
      RECT 653.888 210.096 654.888 211.096 ;
      RECT 653.888 212.096 654.888 213.096 ;
      RECT 653.888 214.096 654.888 215.096 ;
      RECT 653.888 216.096 654.888 217.096 ;
      RECT 651.888 97.676 652.888 98.676 ;
      RECT 651.888 99.676 652.888 100.676 ;
      RECT 651.888 101.676 652.888 102.676 ;
      RECT 651.888 103.676 652.888 104.676 ;
      RECT 651.888 138.5 652.888 139.5 ;
      RECT 651.888 140.5 652.888 141.5 ;
      RECT 651.888 142.5 652.888 143.5 ;
      RECT 651.888 144.5 652.888 145.5 ;
      RECT 651.888 210.096 652.888 211.096 ;
      RECT 651.888 212.096 652.888 213.096 ;
      RECT 651.888 214.096 652.888 215.096 ;
      RECT 651.888 216.096 652.888 217.096 ;
      RECT 576.292 97.676 577.292 98.676 ;
      RECT 576.292 99.676 577.292 100.676 ;
      RECT 576.292 101.676 577.292 102.676 ;
      RECT 576.292 103.676 577.292 104.676 ;
      RECT 574.292 97.676 575.292 98.676 ;
      RECT 574.292 99.676 575.292 100.676 ;
      RECT 574.292 101.676 575.292 102.676 ;
      RECT 574.292 103.676 575.292 104.676 ;
      RECT 572.292 97.676 573.292 98.676 ;
      RECT 572.292 99.676 573.292 100.676 ;
      RECT 572.292 101.676 573.292 102.676 ;
      RECT 572.292 103.676 573.292 104.676 ;
      RECT 570.292 97.676 571.292 98.676 ;
      RECT 570.292 99.676 571.292 100.676 ;
      RECT 570.292 101.676 571.292 102.676 ;
      RECT 570.292 103.676 571.292 104.676 ;
      RECT 555.112 131.676 556.112 132.676 ;
      RECT 555.112 133.676 556.112 134.676 ;
      RECT 555.112 135.676 556.112 136.676 ;
      RECT 555.112 137.676 556.112 138.676 ;
      RECT 553.112 131.676 554.112 132.676 ;
      RECT 553.112 133.676 554.112 134.676 ;
      RECT 553.112 135.676 554.112 136.676 ;
      RECT 553.112 137.676 554.112 138.676 ;
      RECT 551.112 131.676 552.112 132.676 ;
      RECT 551.112 133.676 552.112 134.676 ;
      RECT 551.112 135.676 552.112 136.676 ;
      RECT 551.112 137.676 552.112 138.676 ;
      RECT 549.112 131.676 550.112 132.676 ;
      RECT 549.112 133.676 550.112 134.676 ;
      RECT 549.112 135.676 550.112 136.676 ;
      RECT 549.112 137.676 550.112 138.676 ;
      RECT 358.048 45.5 359.048 46.5 ;
      RECT 358.048 47.5 359.048 48.5 ;
      RECT 358.048 49.5 359.048 50.5 ;
      RECT 358.048 51.5 359.048 52.5 ;
      RECT 356.048 45.5 357.048 46.5 ;
      RECT 356.048 47.5 357.048 48.5 ;
      RECT 356.048 49.5 357.048 50.5 ;
      RECT 356.048 51.5 357.048 52.5 ;
      RECT 354.048 45.5 355.048 46.5 ;
      RECT 354.048 47.5 355.048 48.5 ;
      RECT 354.048 49.5 355.048 50.5 ;
      RECT 354.048 51.5 355.048 52.5 ;
      RECT 352.048 45.5 353.048 46.5 ;
      RECT 352.048 47.5 353.048 48.5 ;
      RECT 352.048 49.5 353.048 50.5 ;
      RECT 352.048 51.5 353.048 52.5 ;
      RECT 335.112 131.676 336.112 132.676 ;
      RECT 335.112 133.676 336.112 134.676 ;
      RECT 335.112 135.676 336.112 136.676 ;
      RECT 335.112 137.676 336.112 138.676 ;
      RECT 333.112 131.676 334.112 132.676 ;
      RECT 333.112 133.676 334.112 134.676 ;
      RECT 333.112 135.676 334.112 136.676 ;
      RECT 333.112 137.676 334.112 138.676 ;
      RECT 331.112 131.676 332.112 132.676 ;
      RECT 331.112 133.676 332.112 134.676 ;
      RECT 331.112 135.676 332.112 136.676 ;
      RECT 331.112 137.676 332.112 138.676 ;
      RECT 329.112 131.676 330.112 132.676 ;
      RECT 329.112 133.676 330.112 134.676 ;
      RECT 329.112 135.676 330.112 136.676 ;
      RECT 329.112 137.676 330.112 138.676 ;
      RECT 137.04 45.5 138.04 46.5 ;
      RECT 137.04 47.5 138.04 48.5 ;
      RECT 137.04 49.5 138.04 50.5 ;
      RECT 137.04 51.5 138.04 52.5 ;
      RECT 135.04 45.5 136.04 46.5 ;
      RECT 135.04 47.5 136.04 48.5 ;
      RECT 135.04 49.5 136.04 50.5 ;
      RECT 135.04 51.5 136.04 52.5 ;
      RECT 133.04 45.5 134.04 46.5 ;
      RECT 133.04 47.5 134.04 48.5 ;
      RECT 133.04 49.5 134.04 50.5 ;
      RECT 133.04 51.5 134.04 52.5 ;
      RECT 131.04 45.5 132.04 46.5 ;
      RECT 131.04 47.5 132.04 48.5 ;
      RECT 131.04 49.5 132.04 50.5 ;
      RECT 131.04 51.5 132.04 52.5 ;
      RECT 115.112 131.676 116.112 132.676 ;
      RECT 115.112 133.676 116.112 134.676 ;
      RECT 115.112 135.676 116.112 136.676 ;
      RECT 115.112 137.676 116.112 138.676 ;
      RECT 113.112 131.676 114.112 132.676 ;
      RECT 113.112 133.676 114.112 134.676 ;
      RECT 113.112 135.676 114.112 136.676 ;
      RECT 113.112 137.676 114.112 138.676 ;
      RECT 111.112 131.676 112.112 132.676 ;
      RECT 111.112 133.676 112.112 134.676 ;
      RECT 111.112 135.676 112.112 136.676 ;
      RECT 111.112 137.676 112.112 138.676 ;
      RECT 109.112 131.676 110.112 132.676 ;
      RECT 109.112 133.676 110.112 134.676 ;
      RECT 109.112 135.676 110.112 136.676 ;
      RECT 109.112 137.676 110.112 138.676 ;
    LAYER Cont ;
      RECT 1206.928 131.676 1207.928 132.676 ;
      RECT 1206.928 133.676 1207.928 134.676 ;
      RECT 1206.928 135.676 1207.928 136.676 ;
      RECT 1206.928 137.676 1207.928 138.676 ;
      RECT 1204.928 131.676 1205.928 132.676 ;
      RECT 1204.928 133.676 1205.928 134.676 ;
      RECT 1204.928 135.676 1205.928 136.676 ;
      RECT 1204.928 137.676 1205.928 138.676 ;
      RECT 1202.928 131.676 1203.928 132.676 ;
      RECT 1202.928 133.676 1203.928 134.676 ;
      RECT 1202.928 135.676 1203.928 136.676 ;
      RECT 1202.928 137.676 1203.928 138.676 ;
      RECT 1200.928 131.676 1201.928 132.676 ;
      RECT 1200.928 133.676 1201.928 134.676 ;
      RECT 1200.928 135.676 1201.928 136.676 ;
      RECT 1200.928 137.676 1201.928 138.676 ;
      RECT 1117.536 46.62 1118.536 47.62 ;
      RECT 1117.536 48.62 1118.536 49.62 ;
      RECT 1117.536 50.62 1118.536 51.62 ;
      RECT 1117.536 52.62 1118.536 53.62 ;
      RECT 1115.536 46.62 1116.536 47.62 ;
      RECT 1115.536 48.62 1116.536 49.62 ;
      RECT 1115.536 50.62 1116.536 51.62 ;
      RECT 1115.536 52.62 1116.536 53.62 ;
      RECT 1113.536 46.62 1114.536 47.62 ;
      RECT 1113.536 48.62 1114.536 49.62 ;
      RECT 1113.536 50.62 1114.536 51.62 ;
      RECT 1113.536 52.62 1114.536 53.62 ;
      RECT 1111.536 46.62 1112.536 47.62 ;
      RECT 1111.536 48.62 1112.536 49.62 ;
      RECT 1111.536 50.62 1112.536 51.62 ;
      RECT 1111.536 52.62 1112.536 53.62 ;
      RECT 986.928 131.676 987.928 132.676 ;
      RECT 986.928 133.676 987.928 134.676 ;
      RECT 986.928 135.676 987.928 136.676 ;
      RECT 986.928 137.676 987.928 138.676 ;
      RECT 984.928 131.676 985.928 132.676 ;
      RECT 984.928 133.676 985.928 134.676 ;
      RECT 984.928 135.676 985.928 136.676 ;
      RECT 984.928 137.676 985.928 138.676 ;
      RECT 982.928 131.676 983.928 132.676 ;
      RECT 982.928 133.676 983.928 134.676 ;
      RECT 982.928 135.676 983.928 136.676 ;
      RECT 982.928 137.676 983.928 138.676 ;
      RECT 980.928 131.676 981.928 132.676 ;
      RECT 980.928 133.676 981.928 134.676 ;
      RECT 980.928 135.676 981.928 136.676 ;
      RECT 980.928 137.676 981.928 138.676 ;
      RECT 905.608 138.4 906.608 139.4 ;
      RECT 905.608 140.4 906.608 141.4 ;
      RECT 905.608 142.4 906.608 143.4 ;
      RECT 905.608 144.4 906.608 145.4 ;
      RECT 903.608 138.4 904.608 139.4 ;
      RECT 903.608 140.4 904.608 141.4 ;
      RECT 903.608 142.4 904.608 143.4 ;
      RECT 903.608 144.4 904.608 145.4 ;
      RECT 901.608 138.4 902.608 139.4 ;
      RECT 901.608 140.4 902.608 141.4 ;
      RECT 901.608 142.4 902.608 143.4 ;
      RECT 901.608 144.4 902.608 145.4 ;
      RECT 899.608 138.4 900.608 139.4 ;
      RECT 899.608 140.4 900.608 141.4 ;
      RECT 899.608 142.4 900.608 143.4 ;
      RECT 899.608 144.4 900.608 145.4 ;
      RECT 787.668 35.676 788.668 36.676 ;
      RECT 787.668 37.676 788.668 38.676 ;
      RECT 787.668 39.676 788.668 40.676 ;
      RECT 787.668 41.676 788.668 42.676 ;
      RECT 785.668 35.676 786.668 36.676 ;
      RECT 785.668 37.676 786.668 38.676 ;
      RECT 785.668 39.676 786.668 40.676 ;
      RECT 785.668 41.676 786.668 42.676 ;
      RECT 783.668 35.676 784.668 36.676 ;
      RECT 783.668 37.676 784.668 38.676 ;
      RECT 783.668 39.676 784.668 40.676 ;
      RECT 783.668 41.676 784.668 42.676 ;
      RECT 781.668 35.676 782.668 36.676 ;
      RECT 781.668 37.676 782.668 38.676 ;
      RECT 781.668 39.676 782.668 40.676 ;
      RECT 781.668 41.676 782.668 42.676 ;
      RECT 769.292 138.4 770.292 139.4 ;
      RECT 769.292 140.4 770.292 141.4 ;
      RECT 769.292 142.4 770.292 143.4 ;
      RECT 769.292 144.4 770.292 145.4 ;
      RECT 767.292 138.4 768.292 139.4 ;
      RECT 767.292 140.4 768.292 141.4 ;
      RECT 767.292 142.4 768.292 143.4 ;
      RECT 767.292 144.4 768.292 145.4 ;
      RECT 765.292 138.4 766.292 139.4 ;
      RECT 765.292 140.4 766.292 141.4 ;
      RECT 765.292 142.4 766.292 143.4 ;
      RECT 765.292 144.4 766.292 145.4 ;
      RECT 763.292 138.4 764.292 139.4 ;
      RECT 763.292 140.4 764.292 141.4 ;
      RECT 763.292 142.4 764.292 143.4 ;
      RECT 763.292 144.4 764.292 145.4 ;
      RECT 707.752 35.676 708.752 36.676 ;
      RECT 707.752 37.676 708.752 38.676 ;
      RECT 707.752 39.676 708.752 40.676 ;
      RECT 707.752 41.676 708.752 42.676 ;
      RECT 705.752 35.676 706.752 36.676 ;
      RECT 705.752 37.676 706.752 38.676 ;
      RECT 705.752 39.676 706.752 40.676 ;
      RECT 705.752 41.676 706.752 42.676 ;
      RECT 703.752 35.676 704.752 36.676 ;
      RECT 703.752 37.676 704.752 38.676 ;
      RECT 703.752 39.676 704.752 40.676 ;
      RECT 703.752 41.676 704.752 42.676 ;
      RECT 701.752 35.676 702.752 36.676 ;
      RECT 701.752 37.676 702.752 38.676 ;
      RECT 701.752 39.676 702.752 40.676 ;
      RECT 701.752 41.676 702.752 42.676 ;
      RECT 688.588 206.772 689.588 207.772 ;
      RECT 688.588 208.772 689.588 209.772 ;
      RECT 688.588 210.772 689.588 211.772 ;
      RECT 688.588 212.772 689.588 213.772 ;
      RECT 686.588 206.772 687.588 207.772 ;
      RECT 686.588 208.772 687.588 209.772 ;
      RECT 686.588 210.772 687.588 211.772 ;
      RECT 686.588 212.772 687.588 213.772 ;
      RECT 685.8 138.5 686.8 139.5 ;
      RECT 685.8 140.5 686.8 141.5 ;
      RECT 685.8 142.5 686.8 143.5 ;
      RECT 685.8 144.5 686.8 145.5 ;
      RECT 684.588 206.772 685.588 207.772 ;
      RECT 684.588 208.772 685.588 209.772 ;
      RECT 684.588 210.772 685.588 211.772 ;
      RECT 684.588 212.772 685.588 213.772 ;
      RECT 683.8 138.5 684.8 139.5 ;
      RECT 683.8 140.5 684.8 141.5 ;
      RECT 683.8 142.5 684.8 143.5 ;
      RECT 683.8 144.5 684.8 145.5 ;
      RECT 682.588 206.772 683.588 207.772 ;
      RECT 682.588 208.772 683.588 209.772 ;
      RECT 682.588 210.772 683.588 211.772 ;
      RECT 682.588 212.772 683.588 213.772 ;
      RECT 681.8 138.5 682.8 139.5 ;
      RECT 681.8 140.5 682.8 141.5 ;
      RECT 681.8 142.5 682.8 143.5 ;
      RECT 681.8 144.5 682.8 145.5 ;
      RECT 679.8 138.5 680.8 139.5 ;
      RECT 679.8 140.5 680.8 141.5 ;
      RECT 679.8 142.5 680.8 143.5 ;
      RECT 679.8 144.5 680.8 145.5 ;
      RECT 648.64 210.096 649.64 211.096 ;
      RECT 648.64 212.096 649.64 213.096 ;
      RECT 648.64 214.096 649.64 215.096 ;
      RECT 648.64 216.096 649.64 217.096 ;
      RECT 646.64 210.096 647.64 211.096 ;
      RECT 646.64 212.096 647.64 213.096 ;
      RECT 646.64 214.096 647.64 215.096 ;
      RECT 646.64 216.096 647.64 217.096 ;
      RECT 644.64 210.096 645.64 211.096 ;
      RECT 644.64 212.096 645.64 213.096 ;
      RECT 644.64 214.096 645.64 215.096 ;
      RECT 644.64 216.096 645.64 217.096 ;
      RECT 642.64 210.096 643.64 211.096 ;
      RECT 642.64 212.096 643.64 213.096 ;
      RECT 642.64 214.096 643.64 215.096 ;
      RECT 642.64 216.096 643.64 217.096 ;
      RECT 566.928 131.676 567.928 132.676 ;
      RECT 566.928 133.676 567.928 134.676 ;
      RECT 566.928 135.676 567.928 136.676 ;
      RECT 566.928 137.676 567.928 138.676 ;
      RECT 564.928 131.676 565.928 132.676 ;
      RECT 564.928 133.676 565.928 134.676 ;
      RECT 564.928 135.676 565.928 136.676 ;
      RECT 564.928 137.676 565.928 138.676 ;
      RECT 562.928 131.676 563.928 132.676 ;
      RECT 562.928 133.676 563.928 134.676 ;
      RECT 562.928 135.676 563.928 136.676 ;
      RECT 562.928 137.676 563.928 138.676 ;
      RECT 560.928 131.676 561.928 132.676 ;
      RECT 560.928 133.676 561.928 134.676 ;
      RECT 560.928 135.676 561.928 136.676 ;
      RECT 560.928 137.676 561.928 138.676 ;
      RECT 528.28 25.536 529.28 26.536 ;
      RECT 528.28 27.536 529.28 28.536 ;
      RECT 528.28 29.536 529.28 30.536 ;
      RECT 528.28 31.536 529.28 32.536 ;
      RECT 526.28 25.536 527.28 26.536 ;
      RECT 526.28 27.536 527.28 28.536 ;
      RECT 526.28 29.536 527.28 30.536 ;
      RECT 526.28 31.536 527.28 32.536 ;
      RECT 524.28 25.536 525.28 26.536 ;
      RECT 524.28 27.536 525.28 28.536 ;
      RECT 524.28 29.536 525.28 30.536 ;
      RECT 524.28 31.536 525.28 32.536 ;
      RECT 522.28 25.536 523.28 26.536 ;
      RECT 522.28 27.536 523.28 28.536 ;
      RECT 522.28 29.536 523.28 30.536 ;
      RECT 522.28 31.536 523.28 32.536 ;
      RECT 370.748 45.5 371.748 46.5 ;
      RECT 370.748 47.5 371.748 48.5 ;
      RECT 370.748 49.5 371.748 50.5 ;
      RECT 370.748 51.5 371.748 52.5 ;
      RECT 368.748 45.5 369.748 46.5 ;
      RECT 368.748 47.5 369.748 48.5 ;
      RECT 368.748 49.5 369.748 50.5 ;
      RECT 368.748 51.5 369.748 52.5 ;
      RECT 366.748 45.5 367.748 46.5 ;
      RECT 366.748 47.5 367.748 48.5 ;
      RECT 366.748 49.5 367.748 50.5 ;
      RECT 366.748 51.5 367.748 52.5 ;
      RECT 364.748 45.5 365.748 46.5 ;
      RECT 364.748 47.5 365.748 48.5 ;
      RECT 364.748 49.5 365.748 50.5 ;
      RECT 364.748 51.5 365.748 52.5 ;
      RECT 346.928 131.676 347.928 132.676 ;
      RECT 346.928 133.676 347.928 134.676 ;
      RECT 346.928 135.676 347.928 136.676 ;
      RECT 346.928 137.676 347.928 138.676 ;
      RECT 344.928 131.676 345.928 132.676 ;
      RECT 344.928 133.676 345.928 134.676 ;
      RECT 344.928 135.676 345.928 136.676 ;
      RECT 344.928 137.676 345.928 138.676 ;
      RECT 342.928 131.676 343.928 132.676 ;
      RECT 342.928 133.676 343.928 134.676 ;
      RECT 342.928 135.676 343.928 136.676 ;
      RECT 342.928 137.676 343.928 138.676 ;
      RECT 340.928 131.676 341.928 132.676 ;
      RECT 340.928 133.676 341.928 134.676 ;
      RECT 340.928 135.676 341.928 136.676 ;
      RECT 340.928 137.676 341.928 138.676 ;
      RECT 267.152 45.612 268.152 46.612 ;
      RECT 267.152 47.612 268.152 48.612 ;
      RECT 267.152 49.612 268.152 50.612 ;
      RECT 267.152 51.612 268.152 52.612 ;
      RECT 265.152 45.612 266.152 46.612 ;
      RECT 265.152 47.612 266.152 48.612 ;
      RECT 265.152 49.612 266.152 50.612 ;
      RECT 265.152 51.612 266.152 52.612 ;
      RECT 263.152 45.612 264.152 46.612 ;
      RECT 263.152 47.612 264.152 48.612 ;
      RECT 263.152 49.612 264.152 50.612 ;
      RECT 263.152 51.612 264.152 52.612 ;
      RECT 261.152 45.612 262.152 46.612 ;
      RECT 261.152 47.612 262.152 48.612 ;
      RECT 261.152 49.612 262.152 50.612 ;
      RECT 261.152 51.612 262.152 52.612 ;
      RECT 149.74 45.5 150.74 46.5 ;
      RECT 149.74 47.5 150.74 48.5 ;
      RECT 149.74 49.5 150.74 50.5 ;
      RECT 149.74 51.5 150.74 52.5 ;
      RECT 147.74 45.5 148.74 46.5 ;
      RECT 147.74 47.5 148.74 48.5 ;
      RECT 147.74 49.5 148.74 50.5 ;
      RECT 147.74 51.5 148.74 52.5 ;
      RECT 145.74 45.5 146.74 46.5 ;
      RECT 145.74 47.5 146.74 48.5 ;
      RECT 145.74 49.5 146.74 50.5 ;
      RECT 145.74 51.5 146.74 52.5 ;
      RECT 143.74 45.5 144.74 46.5 ;
      RECT 143.74 47.5 144.74 48.5 ;
      RECT 143.74 49.5 144.74 50.5 ;
      RECT 143.74 51.5 144.74 52.5 ;
      RECT 126.928 131.676 127.928 132.676 ;
      RECT 126.928 133.676 127.928 134.676 ;
      RECT 126.928 135.676 127.928 136.676 ;
      RECT 126.928 137.676 127.928 138.676 ;
      RECT 124.928 131.676 125.928 132.676 ;
      RECT 124.928 133.676 125.928 134.676 ;
      RECT 124.928 135.676 125.928 136.676 ;
      RECT 124.928 137.676 125.928 138.676 ;
      RECT 122.928 131.676 123.928 132.676 ;
      RECT 122.928 133.676 123.928 134.676 ;
      RECT 122.928 135.676 123.928 136.676 ;
      RECT 122.928 137.676 123.928 138.676 ;
      RECT 120.928 131.676 121.928 132.676 ;
      RECT 120.928 133.676 121.928 134.676 ;
      RECT 120.928 135.676 121.928 136.676 ;
      RECT 120.928 137.676 121.928 138.676 ;
    LAYER Metal1 ;
      RECT 1111.05 25.05 1119.05 54.1 ;
      RECT 521.8 25.05 1119.05 33.05 ;
      RECT 260.65 35.2 268.65 53.1 ;
      RECT 260.65 35.2 789.15 43.2 ;
      RECT 1188.612 131.176 1208.428 139.176 ;
      RECT 968.612 131.176 988.428 139.176 ;
      RECT 762.792 137.9 907.108 145.9 ;
      RECT 670.056 206.272 690.088 214.272 ;
      RECT 651.388 138 687.3 146 ;
      RECT 569.792 97.176 659.388 105.176 ;
      RECT 642.14 209.596 659.388 217.596 ;
      RECT 548.612 131.176 568.428 139.176 ;
      RECT 351.548 45 372.248 53 ;
      RECT 328.612 131.176 348.428 139.176 ;
      RECT 130.54 45 151.24 53 ;
      RECT 108.612 131.176 128.428 139.176 ;
  END
END MoS2DFlipFlop

MACRO MoS2Inverter
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MoS2Inverter 0 0 ;
  SIZE 160 BY 280 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 30 0 40 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 0 160 20 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Contact ;
        RECT 143 211.225 144 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 143 213.225 144 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 143 215.225 144 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 143 217.225 144 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 143 261.65 144 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 143 263.65 144 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 143 265.65 144 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 143 267.65 144 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 141 211.225 142 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 141 213.225 142 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 141 215.225 142 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 141 217.225 142 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 141 261.65 142 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 141 263.65 142 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 141 265.65 142 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 141 267.65 142 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 139 211.225 140 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 139 213.225 140 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 139 215.225 140 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 139 217.225 140 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 139 261.65 140 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 139 263.65 140 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 139 265.65 140 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 139 267.65 140 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 137 211.225 138 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 137 213.225 138 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 137 215.225 138 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 137 217.225 138 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 137 261.65 138 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 137 263.65 138 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 137 265.65 138 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 137 267.65 138 268.65 ;
    END
    PORT
      LAYER NSD ;
        RECT 70 60 80 105.55 ;
    END
    PORT
      LAYER NSD ;
        RECT 70 95.55 145.45 105.55 ;
    END
    PORT
      LAYER NSD ;
        RECT 135.45 95.55 145.45 219.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 260 160 280 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 136.5 210.725 144.5 269.15 ;
    END
  END VDD
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER NSD ;
        RECT 50 39.985 60 90 ;
    END
  END VOUT
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 30 160 40 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 70 160 80 208.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 110 160 120 208.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 30 198.95 120 208.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 230 160 250 ;
    END
  END VSS
  PIN VIN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 39 43.35 51 105 ;
        RECT 19 43.35 51 55.35 ;
        RECT 19 43.35 31 105 ;
    END
  END VIN
  OBS
    LAYER Gate ;
      RECT 79 195 111 205 ;
      RECT 99 145 111 205 ;
      RECT 39 195 71 205 ;
      RECT 59 45 71 205 ;
      RECT 19 145 31 205 ;
      RECT 79 145 91 205 ;
      RECT 39 145 51 205 ;
      RECT 59 145 91 155 ;
      RECT 19 145 51 155 ;
      RECT 25 114.75 71 124.75 ;
      RECT 10 114 20 125 ;
      RECT 136 210 145 220 ;
      RECT 136 260 145 270 ;
    LAYER NSD ;
      RECT 90 142.25 100 190 ;
      RECT 50 142.25 60 190 ;
      RECT 10 60 20 190 ;
      RECT 10 142.25 100 152.25 ;
      RECT 24 114 35 125 ;
    LAYER Contact ;
      RECT 18.5 115.265 19.5 116.265 ;
      RECT 18.5 117.265 19.5 118.265 ;
      RECT 18.5 119.265 19.5 120.265 ;
      RECT 18.5 121.265 19.5 122.265 ;
      RECT 18.5 123.265 19.5 124.265 ;
      RECT 16.5 115.265 17.5 116.265 ;
      RECT 16.5 117.265 17.5 118.265 ;
      RECT 16.5 119.265 17.5 120.265 ;
      RECT 16.5 121.265 17.5 122.265 ;
      RECT 16.5 123.265 17.5 124.265 ;
      RECT 14.5 115.265 15.5 116.265 ;
      RECT 14.5 117.265 15.5 118.265 ;
      RECT 14.5 119.265 15.5 120.265 ;
      RECT 14.5 121.265 15.5 122.265 ;
      RECT 14.5 123.265 15.5 124.265 ;
      RECT 12.5 115.265 13.5 116.265 ;
      RECT 12.5 117.265 13.5 118.265 ;
      RECT 12.5 119.265 13.5 120.265 ;
      RECT 12.5 121.265 13.5 122.265 ;
      RECT 12.5 123.265 13.5 124.265 ;
      RECT 10.5 115.265 11.5 116.265 ;
      RECT 10.5 117.265 11.5 118.265 ;
      RECT 10.5 119.265 11.5 120.265 ;
      RECT 10.5 121.265 11.5 122.265 ;
      RECT 10.5 123.265 11.5 124.265 ;
      RECT 79 195 111 205 ;
      RECT 99 145 111 205 ;
      RECT 39 195 71 205 ;
      RECT 59 45 71 205 ;
      RECT 19 145 31 205 ;
      RECT 79 145 91 205 ;
      RECT 39 145 51 205 ;
      RECT 59 145 91 155 ;
      RECT 19 145 51 155 ;
      RECT 25 114.75 71 124.75 ;
        RECT 39 43.35 51 105 ;
        RECT 19 43.35 51 55.35 ;
        RECT 19 43.35 31 105 ;
    LAYER Cont ;
      RECT 33.5 115.265 34.5 116.265 ;
      RECT 33.5 117.265 34.5 118.265 ;
      RECT 33.5 119.265 34.5 120.265 ;
      RECT 33.5 121.265 34.5 122.265 ;
      RECT 33.5 123.265 34.5 124.265 ;
      RECT 31.5 115.265 32.5 116.265 ;
      RECT 31.5 117.265 32.5 118.265 ;
      RECT 31.5 119.265 32.5 120.265 ;
      RECT 31.5 121.265 32.5 122.265 ;
      RECT 31.5 123.265 32.5 124.265 ;
      RECT 29.5 115.265 30.5 116.265 ;
      RECT 29.5 117.265 30.5 118.265 ;
      RECT 29.5 119.265 30.5 120.265 ;
      RECT 29.5 121.265 30.5 122.265 ;
      RECT 29.5 123.265 30.5 124.265 ;
      RECT 27.5 115.265 28.5 116.265 ;
      RECT 27.5 117.265 28.5 118.265 ;
      RECT 27.5 119.265 28.5 120.265 ;
      RECT 27.5 121.265 28.5 122.265 ;
      RECT 27.5 123.265 28.5 124.265 ;
      RECT 25.5 115.265 26.5 116.265 ;
      RECT 25.5 117.265 26.5 118.265 ;
      RECT 25.5 119.265 26.5 120.265 ;
      RECT 25.5 121.265 26.5 122.265 ;
      RECT 25.5 123.265 26.5 124.265 ;
      RECT 90 142.25 100 190 ;
      RECT 50 142.25 60 190 ;
      RECT 10 60 20 190 ;
      RECT 10 142.25 100 152.25 ;
        RECT 30 0 40 90 ;
        RECT 0 0 160 20 ;
        RECT 70 60 80 105.55 ;
        RECT 70 95.55 145.45 105.55 ;
        RECT 135.45 95.55 145.45 219.1 ;
        RECT 0 260 160 280 ;
        RECT 50 39.985 60 90 ;
        RECT 30 160 40 250 ;
        RECT 70 160 80 208.95 ;
        RECT 110 160 120 208.95 ;
        RECT 30 198.95 120 208.95 ;
        RECT 0 230 160 250 ;
    LAYER Metal1 ;
      RECT 10 114.765 35 124.765 ;
  END
END MoS2Inverter

MACRO MoS2Nand
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MoS2Nand 0 0 ;
  SIZE 220 BY 280 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 10 0 20 190 ;
    END
    PORT
      LAYER NSD ;
        RECT 50 0 60 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 0 220 20 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Contact ;
        RECT 184.355 212.915 185.355 213.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 184.355 214.915 185.355 215.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 184.355 216.915 185.355 217.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 184.355 218.915 185.355 219.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 184.355 261.91 185.355 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 184.355 263.91 185.355 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 184.355 265.91 185.355 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 184.355 267.91 185.355 268.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 182.355 212.915 183.355 213.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 182.355 214.915 183.355 215.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 182.355 216.915 183.355 217.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 182.355 218.915 183.355 219.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 182.355 261.91 183.355 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 182.355 263.91 183.355 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 182.355 265.91 183.355 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 182.355 267.91 183.355 268.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 180.355 212.915 181.355 213.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 180.355 214.915 181.355 215.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 180.355 216.915 181.355 217.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 180.355 218.915 181.355 219.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 180.355 261.91 181.355 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 180.355 263.91 181.355 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 180.355 265.91 181.355 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 180.355 267.91 181.355 268.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 178.355 212.915 179.355 213.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 178.355 214.915 179.355 215.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 178.355 216.915 179.355 217.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 178.355 218.915 179.355 219.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 178.355 261.91 179.355 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 178.355 263.91 179.355 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 178.355 265.91 179.355 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 178.355 267.91 179.355 268.91 ;
    END
    PORT
      LAYER NSD ;
        RECT 150 60 160 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 150 98.9 186.85 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 176.85 98.9 186.85 220.75 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 260 220 280 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 177.855 212.415 185.855 269.41 ;
    END
  END VDD
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6 LAYER NSD ;
    PORT
      LAYER NSD ;
        RECT 90 96.35 140 106.35 ;
        RECT 130 60 140 106.35 ;
        RECT 90 60 100 106.35 ;
    END
  END VOUT
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 70 160 80 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 110 160 120 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 150 160 160 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 70 198.1 160 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 230 220 250 ;
    END
  END VSS
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 99 45 111 105 ;
        RECT 79 45 111 55 ;
        RECT 39 122 91 134 ;
        RECT 79 45 91 134 ;
        RECT 39 122 51 205 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 39 45 51 105 ;
        RECT 19 45 51 55 ;
        RECT 19 45 31 205 ;
    END
  END B
  OBS
    LAYER Gate ;
      RECT 119 195 151 205 ;
      RECT 139 145 151 205 ;
      RECT 79 195 111 205 ;
      RECT 99 145 111 205 ;
      RECT 59 145 71 205 ;
      RECT 119 122.6 131 205 ;
      RECT 79 145 91 205 ;
      RECT 99 145 131 155 ;
      RECT 59 145 91 155 ;
      RECT 119 122.6 151 134.6 ;
      RECT 139 45 151 134.6 ;
      RECT 108 131 117 140 ;
      RECT 40 207 49 216 ;
      RECT 31 33 40 42 ;
      RECT 177 212 186 221 ;
      RECT 177 260 186 270 ;
    LAYER NSD ;
      RECT 130 141.75 140 190 ;
      RECT 90 141.75 100 190 ;
      RECT 50 141.75 60 190 ;
      RECT 50 141.75 140 151.75 ;
      RECT 108.6 131.2 116.6 151.75 ;
      RECT 30 96.35 80 106.35 ;
      RECT 70 42.05 80 106.35 ;
      RECT 30 60 40 106.35 ;
      RECT 110 42.05 120 90 ;
      RECT 70 42.05 120 52.05 ;
      RECT 30 160 40 190 ;
      RECT 120 131 128 139 ;
      RECT 40 196 49 205 ;
      RECT 31 44 40 55 ;
      RECT 119 131 129 140 ;
    LAYER Contact ;
      RECT 115.11 131.675 116.11 132.675 ;
      RECT 115.11 133.675 116.11 134.675 ;
      RECT 115.11 135.675 116.11 136.675 ;
      RECT 115.11 137.675 116.11 138.675 ;
      RECT 113.11 131.675 114.11 132.675 ;
      RECT 113.11 133.675 114.11 134.675 ;
      RECT 113.11 135.675 114.11 136.675 ;
      RECT 113.11 137.675 114.11 138.675 ;
      RECT 111.11 131.675 112.11 132.675 ;
      RECT 111.11 133.675 112.11 134.675 ;
      RECT 111.11 135.675 112.11 136.675 ;
      RECT 111.11 137.675 112.11 138.675 ;
      RECT 109.11 131.675 110.11 132.675 ;
      RECT 109.11 133.675 110.11 134.675 ;
      RECT 109.11 135.675 110.11 136.675 ;
      RECT 109.11 137.675 110.11 138.675 ;
      RECT 119 195 151 205 ;
      RECT 139 145 151 205 ;
      RECT 79 195 111 205 ;
      RECT 99 145 111 205 ;
      RECT 59 145 71 205 ;
      RECT 119 122.6 131 205 ;
      RECT 79 145 91 205 ;
      RECT 99 145 131 155 ;
      RECT 59 145 91 155 ;
      RECT 119 122.6 151 134.6 ;
      RECT 139 45 151 134.6 ;
        RECT 99 45 111 105 ;
        RECT 79 45 111 55 ;
        RECT 39 122 91 134 ;
        RECT 79 45 91 134 ;
        RECT 39 122 51 205 ;
        RECT 39 45 51 105 ;
        RECT 19 45 51 55 ;
        RECT 19 45 31 205 ;
    LAYER Cont ;
      RECT 126.925 131.675 127.925 132.675 ;
      RECT 126.925 133.675 127.925 134.675 ;
      RECT 126.925 135.675 127.925 136.675 ;
      RECT 126.925 137.675 127.925 138.675 ;
      RECT 124.925 131.675 125.925 132.675 ;
      RECT 124.925 133.675 125.925 134.675 ;
      RECT 124.925 135.675 125.925 136.675 ;
      RECT 124.925 137.675 125.925 138.675 ;
      RECT 122.925 131.675 123.925 132.675 ;
      RECT 122.925 133.675 123.925 134.675 ;
      RECT 122.925 135.675 123.925 136.675 ;
      RECT 122.925 137.675 123.925 138.675 ;
      RECT 120.925 131.675 121.925 132.675 ;
      RECT 120.925 133.675 121.925 134.675 ;
      RECT 120.925 135.675 121.925 136.675 ;
      RECT 120.925 137.675 121.925 138.675 ;
      RECT 130 141.75 140 190 ;
      RECT 90 141.75 100 190 ;
      RECT 50 141.75 60 190 ;
      RECT 50 141.75 140 151.75 ;
      RECT 108.6 131.2 116.6 151.75 ;
      RECT 30 96.35 80 106.35 ;
      RECT 70 42.05 80 106.35 ;
      RECT 30 60 40 106.35 ;
      RECT 110 42.05 120 90 ;
      RECT 70 42.05 120 52.05 ;
      RECT 30 160 40 190 ;
      RECT 120 131 128 139 ;
      RECT 10 0 20 190 ;
        RECT 50 0 60 90 ;
        RECT 0 0 220 20 ;
        RECT 150 60 160 108.9 ;
        RECT 150 98.9 186.85 108.9 ;
        RECT 176.85 98.9 186.85 220.75 ;
        RECT 0 260 220 280 ;
        RECT 90 96.35 140 106.35 ;
        RECT 130 60 140 106.35 ;
        RECT 90 60 100 106.35 ;
        RECT 70 160 80 250 ;
        RECT 110 160 120 208.1 ;
        RECT 150 160 160 208.1 ;
        RECT 70 198.1 160 208.1 ;
        RECT 0 230 220 250 ;
    LAYER Metal1 ;
      RECT 108.61 131.175 128.425 139.175 ;
  END
END MoS2Nand

MACRO MoS2Nor
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MoS2Nor 0 0 ;
  SIZE 220 BY 280 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 19 100.5 71 112.5 ;
        RECT 59 45 71 112.5 ;
        RECT 19 45 31 112.5 ;
      LAYER Metal1 ;
        RECT 9.425 102.965 28.01 110.965 ;
      LAYER NSD ;
        RECT 9.425 102.965 17.425 110.965 ;
      LAYER Cont ;
        RECT 20.51 109.465 21.51 110.465 ;
        RECT 20.51 107.465 21.51 108.465 ;
        RECT 20.51 105.465 21.51 106.465 ;
        RECT 20.51 103.465 21.51 104.465 ;
        RECT 22.51 109.465 23.51 110.465 ;
        RECT 22.51 107.465 23.51 108.465 ;
        RECT 22.51 105.465 23.51 106.465 ;
        RECT 22.51 103.465 23.51 104.465 ;
        RECT 24.51 109.465 25.51 110.465 ;
        RECT 24.51 107.465 25.51 108.465 ;
        RECT 24.51 105.465 25.51 106.465 ;
        RECT 24.51 103.465 25.51 104.465 ;
        RECT 26.51 109.465 27.51 110.465 ;
        RECT 26.51 107.465 27.51 108.465 ;
        RECT 26.51 105.465 27.51 106.465 ;
        RECT 26.51 103.465 27.51 104.465 ;
      LAYER Contact ;
        RECT 9.925 109.465 10.925 110.465 ;
        RECT 9.925 107.465 10.925 108.465 ;
        RECT 9.925 105.465 10.925 106.465 ;
        RECT 9.925 103.465 10.925 104.465 ;
        RECT 11.925 109.465 12.925 110.465 ;
        RECT 11.925 107.465 12.925 108.465 ;
        RECT 11.925 105.465 12.925 106.465 ;
        RECT 11.925 103.465 12.925 104.465 ;
        RECT 13.925 109.465 14.925 110.465 ;
        RECT 13.925 107.465 14.925 108.465 ;
        RECT 13.925 105.465 14.925 106.465 ;
        RECT 13.925 103.465 14.925 104.465 ;
        RECT 15.925 109.465 16.925 110.465 ;
        RECT 15.925 107.465 16.925 108.465 ;
        RECT 15.925 105.465 16.925 106.465 ;
        RECT 15.925 103.465 16.925 104.465 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 79 27.35 91 105 ;
        RECT 39 27.35 91 39.35 ;
        RECT 39 27.35 51 95.55 ;
      LAYER Metal1 ;
        RECT 28.245 28.835 48.225 36.835 ;
      LAYER NSD ;
        RECT 28.245 28.835 36.245 36.835 ;
      LAYER Cont ;
        RECT 40.725 35.335 41.725 36.335 ;
        RECT 40.725 33.335 41.725 34.335 ;
        RECT 40.725 31.335 41.725 32.335 ;
        RECT 40.725 29.335 41.725 30.335 ;
        RECT 42.725 35.335 43.725 36.335 ;
        RECT 42.725 33.335 43.725 34.335 ;
        RECT 42.725 31.335 43.725 32.335 ;
        RECT 42.725 29.335 43.725 30.335 ;
        RECT 44.725 35.335 45.725 36.335 ;
        RECT 44.725 33.335 45.725 34.335 ;
        RECT 44.725 31.335 45.725 32.335 ;
        RECT 44.725 29.335 45.725 30.335 ;
        RECT 46.725 35.335 47.725 36.335 ;
        RECT 46.725 33.335 47.725 34.335 ;
        RECT 46.725 31.335 47.725 32.335 ;
        RECT 46.725 29.335 47.725 30.335 ;
      LAYER Contact ;
        RECT 28.745 35.335 29.745 36.335 ;
        RECT 28.745 33.335 29.745 34.335 ;
        RECT 28.745 31.335 29.745 32.335 ;
        RECT 28.745 29.335 29.745 30.335 ;
        RECT 30.745 35.335 31.745 36.335 ;
        RECT 30.745 33.335 31.745 34.335 ;
        RECT 30.745 31.335 31.745 32.335 ;
        RECT 30.745 29.335 31.745 30.335 ;
        RECT 32.745 35.335 33.745 36.335 ;
        RECT 32.745 33.335 33.745 34.335 ;
        RECT 32.745 31.335 33.745 32.335 ;
        RECT 32.745 29.335 33.745 30.335 ;
        RECT 34.745 35.335 35.745 36.335 ;
        RECT 34.745 33.335 35.745 34.335 ;
        RECT 34.745 31.335 35.745 32.335 ;
        RECT 34.745 29.335 35.745 30.335 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 10 0 20 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 50 0 60 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 90 0 100 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 0 220 20 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Contact ;
        RECT 147.445 216.875 148.445 217.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 147.445 218.875 148.445 219.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 147.445 220.875 148.445 221.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 147.445 222.875 148.445 223.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 147.445 262.575 148.445 263.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 147.445 264.575 148.445 265.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 147.445 266.575 148.445 267.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 147.445 268.575 148.445 269.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 216.875 146.445 217.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 218.875 146.445 219.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 220.875 146.445 221.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 222.875 146.445 223.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 262.575 146.445 263.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 264.575 146.445 265.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 266.575 146.445 267.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 268.575 146.445 269.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 216.875 144.445 217.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 218.875 144.445 219.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 220.875 144.445 221.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 222.875 144.445 223.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 262.575 144.445 263.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 264.575 144.445 265.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 266.575 144.445 267.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 268.575 144.445 269.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 216.875 142.445 217.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 218.875 142.445 219.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 220.875 142.445 221.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 222.875 142.445 223.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 262.575 142.445 263.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 264.575 142.445 265.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 266.575 142.445 267.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 268.575 142.445 269.575 ;
    END
    PORT
      LAYER NSD ;
        RECT 140 160 150 225.2 ;
    END
    PORT
      LAYER NSD ;
        RECT 180 160 190 207.5 ;
    END
    PORT
      LAYER NSD ;
        RECT 140 197.5 190 207.5 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 260 220 280 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 140.945 216.375 148.945 270.075 ;
    END
  END VDD
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER NSD ;
        RECT 160 112.9 170 190 ;
        RECT 70 112.9 170 122.9 ;
        RECT 70 60 80 122.9 ;
    END
  END VOUT
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 30 160 40 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 70 160 80 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 110 160 120 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 230 220 250 ;
    END
  END VSS
  OBS
    LAYER Gate ;
      RECT 169 145 181 205 ;
      RECT 79 195 161 205 ;
      RECT 149 145 161 205 ;
      RECT 39 195 71 205 ;
      RECT 59 145 71 205 ;
      RECT 19 145 31 205 ;
      RECT 99 193 161 205 ;
      RECT 79 145 91 205 ;
      RECT 39 145 51 205 ;
      RECT 99 145 111 205 ;
      RECT 149 145 181 155 ;
      RECT 59 145 91 155 ;
      RECT 19 145 51 155 ;
    LAYER NSD ;
      RECT 90 134.45 100 190 ;
      RECT 50 134.45 60 190 ;
      RECT 10 134.45 20 190 ;
      RECT 10 134.45 100 144.45 ;
      RECT 30 60 40 144.45 ;
    LAYER Contact ;
      RECT 16.575 145.655 17.575 146.655 ;
      RECT 16.575 147.655 17.575 148.655 ;
      RECT 16.575 149.655 17.575 150.655 ;
      RECT 16.575 151.655 17.575 152.655 ;
      RECT 14.575 145.655 15.575 146.655 ;
      RECT 14.575 147.655 15.575 148.655 ;
      RECT 14.575 149.655 15.575 150.655 ;
      RECT 14.575 151.655 15.575 152.655 ;
      RECT 12.575 145.655 13.575 146.655 ;
      RECT 12.575 147.655 13.575 148.655 ;
      RECT 12.575 149.655 13.575 150.655 ;
      RECT 12.575 151.655 13.575 152.655 ;
      RECT 10.575 145.655 11.575 146.655 ;
      RECT 10.575 147.655 11.575 148.655 ;
      RECT 10.575 149.655 11.575 150.655 ;
      RECT 10.575 151.655 11.575 152.655 ;
    LAYER Cont ;
      RECT 27.52 145.655 28.52 146.655 ;
      RECT 27.52 147.655 28.52 148.655 ;
      RECT 27.52 149.655 28.52 150.655 ;
      RECT 27.52 151.655 28.52 152.655 ;
      RECT 25.52 145.655 26.52 146.655 ;
      RECT 25.52 147.655 26.52 148.655 ;
      RECT 25.52 149.655 26.52 150.655 ;
      RECT 25.52 151.655 26.52 152.655 ;
      RECT 23.52 145.655 24.52 146.655 ;
      RECT 23.52 147.655 24.52 148.655 ;
      RECT 23.52 149.655 24.52 150.655 ;
      RECT 23.52 151.655 24.52 152.655 ;
      RECT 21.52 145.655 22.52 146.655 ;
      RECT 21.52 147.655 22.52 148.655 ;
      RECT 21.52 149.655 22.52 150.655 ;
      RECT 21.52 151.655 22.52 152.655 ;
    LAYER Metal1 ;
      RECT 10.075 145.155 29.02 153.155 ;
  END
END MoS2Nor

MACRO MoS2Or
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MoS2Or 0 0 ;
  SIZE 350 BY 280 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 10 0 20 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 50 0 60 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 90 0 100 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 220 0 230 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 0 350 20 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Contact ;
        RECT 328.2 211.225 329.2 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 328.2 213.225 329.2 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 328.2 215.225 329.2 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 328.2 217.225 329.2 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 328.2 261.65 329.2 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 328.2 263.65 329.2 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 328.2 265.65 329.2 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 328.2 267.65 329.2 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 326.2 211.225 327.2 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 326.2 213.225 327.2 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 326.2 215.225 327.2 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 326.2 217.225 327.2 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 326.2 261.65 327.2 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 326.2 263.65 327.2 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 326.2 265.65 327.2 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 326.2 267.65 327.2 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 324.2 211.225 325.2 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 324.2 213.225 325.2 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 324.2 215.225 325.2 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 324.2 217.225 325.2 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 324.2 261.65 325.2 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 324.2 263.65 325.2 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 324.2 265.65 325.2 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 324.2 267.65 325.2 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 322.2 211.225 323.2 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 322.2 213.225 323.2 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 322.2 215.225 323.2 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 322.2 217.225 323.2 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 322.2 261.65 323.2 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 322.2 263.65 323.2 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 322.2 265.65 323.2 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 322.2 267.65 323.2 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 147.445 216.875 148.445 217.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 147.445 218.875 148.445 219.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 147.445 220.875 148.445 221.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 147.445 222.875 148.445 223.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 147.445 262.575 148.445 263.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 147.445 264.575 148.445 265.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 147.445 266.575 148.445 267.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 147.445 268.575 148.445 269.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 216.875 146.445 217.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 218.875 146.445 219.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 220.875 146.445 221.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 222.875 146.445 223.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 262.575 146.445 263.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 264.575 146.445 265.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 266.575 146.445 267.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 145.445 268.575 146.445 269.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 216.875 144.445 217.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 218.875 144.445 219.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 220.875 144.445 221.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 222.875 144.445 223.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 262.575 144.445 263.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 264.575 144.445 265.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 266.575 144.445 267.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 143.445 268.575 144.445 269.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 216.875 142.445 217.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 218.875 142.445 219.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 220.875 142.445 221.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 222.875 142.445 223.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 262.575 142.445 263.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 264.575 142.445 265.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 266.575 142.445 267.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 141.445 268.575 142.445 269.575 ;
    END
    PORT
      LAYER NSD ;
        RECT 140 160 150 225.2 ;
    END
    PORT
      LAYER NSD ;
        RECT 180 160 190 207.5 ;
    END
    PORT
      LAYER NSD ;
        RECT 140 197.5 190 207.5 ;
    END
    PORT
      LAYER NSD ;
        RECT 260 60 270 105.55 ;
    END
    PORT
      LAYER NSD ;
        RECT 260 95.55 330.55 105.55 ;
    END
    PORT
      LAYER NSD ;
        RECT 320.55 95.55 330.55 219.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 260 350 280 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 140.945 216.375 148.945 270.075 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 321.7 210.725 329.7 269.15 ;
    END
  END VDD
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER NSD ;
        RECT 240 42.165 250 90 ;
    END
  END VOUT
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 30 160 40 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 70 160 80 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 110 160 120 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 220 160 230 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 260 160 270 208.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 300 160 310 208.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 220 198.95 310 208.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 230 350 250 ;
    END
  END VSS
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 19 100.5 71 112.5 ;
        RECT 59 45 71 112.5 ;
        RECT 19 45 31 112.5 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 79 27.35 91 105 ;
        RECT 39 27.35 91 39.35 ;
        RECT 39 27.35 51 95.55 ;
    END
  END B
  OBS
    LAYER Gate ;
      RECT 269 195 301 205 ;
      RECT 289 145 301 205 ;
      RECT 229 195 261 205 ;
      RECT 249 45 261 205 ;
      RECT 209 145 221 205 ;
      RECT 269 145 281 205 ;
      RECT 229 145 241 205 ;
      RECT 249 145 281 155 ;
      RECT 209 145 241 155 ;
      RECT 215 114.75 261 124.75 ;
      RECT 229 43.35 241 105 ;
      RECT 209 43.35 221 105 ;
      RECT 209 43.35 241 55.35 ;
      RECT 169 145 181 205 ;
      RECT 79 195 161 205 ;
      RECT 149 145 161 205 ;
      RECT 39 195 71 205 ;
      RECT 59 145 71 205 ;
      RECT 19 145 31 205 ;
      RECT 99 193 161 205 ;
      RECT 79 145 91 205 ;
      RECT 39 145 51 205 ;
      RECT 99 145 111 205 ;
      RECT 149 145 181 155 ;
      RECT 59 145 91 155 ;
      RECT 19 145 51 155 ;
      RECT 200 114 210 125 ;
      RECT 193 43 204 54 ;
      RECT 10 145 19 153 ;
      RECT 140 262 149 270 ;
      RECT 140 216 149 225 ;
      RECT 321 210 330 219 ;
      RECT 321 261 330 270 ;
    LAYER NSD ;
      RECT 280 142.25 290 190 ;
      RECT 240 142.25 250 190 ;
      RECT 200 60 210 190 ;
      RECT 200 142.25 290 152.25 ;
      RECT 160 43.35 170 190 ;
      RECT 70 112.9 170 122.9 ;
      RECT 70 60 80 122.9 ;
      RECT 160 43.35 203.6 53.35 ;
      RECT 90 134.45 100 190 ;
      RECT 50 134.45 60 190 ;
      RECT 10 134.45 20 190 ;
      RECT 10 134.45 100 144.45 ;
      RECT 30 60 40 144.45 ;
      RECT 215 115 225 125 ;
      RECT 209 43 219 53 ;
      RECT 21 145 29 153 ;
      RECT 20 145 30 154 ;
      RECT 214 114 224 124 ;
      RECT 208 43 218 53 ;
    LAYER Contact ;
      RECT 208.5 115.265 209.5 116.265 ;
      RECT 208.5 117.265 209.5 118.265 ;
      RECT 208.5 119.265 209.5 120.265 ;
      RECT 208.5 121.265 209.5 122.265 ;
      RECT 208.5 123.265 209.5 124.265 ;
      RECT 206.5 115.265 207.5 116.265 ;
      RECT 206.5 117.265 207.5 118.265 ;
      RECT 206.5 119.265 207.5 120.265 ;
      RECT 206.5 121.265 207.5 122.265 ;
      RECT 206.5 123.265 207.5 124.265 ;
      RECT 204.5 115.265 205.5 116.265 ;
      RECT 204.5 117.265 205.5 118.265 ;
      RECT 204.5 119.265 205.5 120.265 ;
      RECT 204.5 121.265 205.5 122.265 ;
      RECT 204.5 123.265 205.5 124.265 ;
      RECT 202.5 115.265 203.5 116.265 ;
      RECT 202.5 117.265 203.5 118.265 ;
      RECT 202.5 119.265 203.5 120.265 ;
      RECT 202.5 121.265 203.5 122.265 ;
      RECT 202.5 123.265 203.5 124.265 ;
      RECT 202.09 43.835 203.09 44.835 ;
      RECT 202.09 45.835 203.09 46.835 ;
      RECT 202.09 47.835 203.09 48.835 ;
      RECT 202.09 49.835 203.09 50.835 ;
      RECT 202.09 51.835 203.09 52.835 ;
      RECT 200.5 115.265 201.5 116.265 ;
      RECT 200.5 117.265 201.5 118.265 ;
      RECT 200.5 119.265 201.5 120.265 ;
      RECT 200.5 121.265 201.5 122.265 ;
      RECT 200.5 123.265 201.5 124.265 ;
      RECT 200.09 43.835 201.09 44.835 ;
      RECT 200.09 45.835 201.09 46.835 ;
      RECT 200.09 47.835 201.09 48.835 ;
      RECT 200.09 49.835 201.09 50.835 ;
      RECT 200.09 51.835 201.09 52.835 ;
      RECT 198.09 43.835 199.09 44.835 ;
      RECT 198.09 45.835 199.09 46.835 ;
      RECT 198.09 47.835 199.09 48.835 ;
      RECT 198.09 49.835 199.09 50.835 ;
      RECT 198.09 51.835 199.09 52.835 ;
      RECT 196.09 43.835 197.09 44.835 ;
      RECT 196.09 45.835 197.09 46.835 ;
      RECT 196.09 47.835 197.09 48.835 ;
      RECT 196.09 49.835 197.09 50.835 ;
      RECT 196.09 51.835 197.09 52.835 ;
      RECT 194.09 43.835 195.09 44.835 ;
      RECT 194.09 45.835 195.09 46.835 ;
      RECT 194.09 47.835 195.09 48.835 ;
      RECT 194.09 49.835 195.09 50.835 ;
      RECT 194.09 51.835 195.09 52.835 ;
      RECT 16.575 145.655 17.575 146.655 ;
      RECT 16.575 147.655 17.575 148.655 ;
      RECT 16.575 149.655 17.575 150.655 ;
      RECT 16.575 151.655 17.575 152.655 ;
      RECT 14.575 145.655 15.575 146.655 ;
      RECT 14.575 147.655 15.575 148.655 ;
      RECT 14.575 149.655 15.575 150.655 ;
      RECT 14.575 151.655 15.575 152.655 ;
      RECT 12.575 145.655 13.575 146.655 ;
      RECT 12.575 147.655 13.575 148.655 ;
      RECT 12.575 149.655 13.575 150.655 ;
      RECT 12.575 151.655 13.575 152.655 ;
      RECT 10.575 145.655 11.575 146.655 ;
      RECT 10.575 147.655 11.575 148.655 ;
      RECT 10.575 149.655 11.575 150.655 ;
      RECT 10.575 151.655 11.575 152.655 ;
      RECT 269 195 301 205 ;
      RECT 289 145 301 205 ;
      RECT 229 195 261 205 ;
      RECT 249 45 261 205 ;
      RECT 209 145 221 205 ;
      RECT 269 145 281 205 ;
      RECT 229 145 241 205 ;
      RECT 249 145 281 155 ;
      RECT 209 145 241 155 ;
      RECT 215 114.75 261 124.75 ;
      RECT 229 43.35 241 105 ;
      RECT 209 43.35 221 105 ;
      RECT 209 43.35 241 55.35 ;
      RECT 169 145 181 205 ;
      RECT 79 195 161 205 ;
      RECT 149 145 161 205 ;
      RECT 39 195 71 205 ;
      RECT 59 145 71 205 ;
      RECT 19 145 31 205 ;
      RECT 99 193 161 205 ;
      RECT 79 145 91 205 ;
      RECT 39 145 51 205 ;
      RECT 99 145 111 205 ;
      RECT 149 145 181 155 ;
      RECT 59 145 91 155 ;
      RECT 19 145 51 155 ;
        RECT 19 100.5 71 112.5 ;
        RECT 59 45 71 112.5 ;
        RECT 19 45 31 112.5 ;
        RECT 79 27.35 91 105 ;
        RECT 39 27.35 91 39.35 ;
        RECT 39 27.35 51 95.55 ;
    LAYER Cont ;
      RECT 223.5 115.265 224.5 116.265 ;
      RECT 223.5 117.265 224.5 118.265 ;
      RECT 223.5 119.265 224.5 120.265 ;
      RECT 223.5 121.265 224.5 122.265 ;
      RECT 223.5 123.265 224.5 124.265 ;
      RECT 221.5 115.265 222.5 116.265 ;
      RECT 221.5 117.265 222.5 118.265 ;
      RECT 221.5 119.265 222.5 120.265 ;
      RECT 221.5 121.265 222.5 122.265 ;
      RECT 221.5 123.265 222.5 124.265 ;
      RECT 219.5 115.265 220.5 116.265 ;
      RECT 219.5 117.265 220.5 118.265 ;
      RECT 219.5 119.265 220.5 120.265 ;
      RECT 219.5 121.265 220.5 122.265 ;
      RECT 219.5 123.265 220.5 124.265 ;
      RECT 217.5 43.835 218.5 44.835 ;
      RECT 217.5 45.835 218.5 46.835 ;
      RECT 217.5 47.835 218.5 48.835 ;
      RECT 217.5 49.835 218.5 50.835 ;
      RECT 217.5 51.835 218.5 52.835 ;
      RECT 217.5 115.265 218.5 116.265 ;
      RECT 217.5 117.265 218.5 118.265 ;
      RECT 217.5 119.265 218.5 120.265 ;
      RECT 217.5 121.265 218.5 122.265 ;
      RECT 217.5 123.265 218.5 124.265 ;
      RECT 215.5 43.835 216.5 44.835 ;
      RECT 215.5 45.835 216.5 46.835 ;
      RECT 215.5 47.835 216.5 48.835 ;
      RECT 215.5 49.835 216.5 50.835 ;
      RECT 215.5 51.835 216.5 52.835 ;
      RECT 215.5 115.265 216.5 116.265 ;
      RECT 215.5 117.265 216.5 118.265 ;
      RECT 215.5 119.265 216.5 120.265 ;
      RECT 215.5 121.265 216.5 122.265 ;
      RECT 215.5 123.265 216.5 124.265 ;
      RECT 213.5 43.835 214.5 44.835 ;
      RECT 213.5 45.835 214.5 46.835 ;
      RECT 213.5 47.835 214.5 48.835 ;
      RECT 213.5 49.835 214.5 50.835 ;
      RECT 213.5 51.835 214.5 52.835 ;
      RECT 211.5 43.835 212.5 44.835 ;
      RECT 211.5 45.835 212.5 46.835 ;
      RECT 211.5 47.835 212.5 48.835 ;
      RECT 211.5 49.835 212.5 50.835 ;
      RECT 211.5 51.835 212.5 52.835 ;
      RECT 209.5 43.835 210.5 44.835 ;
      RECT 209.5 45.835 210.5 46.835 ;
      RECT 209.5 47.835 210.5 48.835 ;
      RECT 209.5 49.835 210.5 50.835 ;
      RECT 209.5 51.835 210.5 52.835 ;
      RECT 27.52 145.655 28.52 146.655 ;
      RECT 27.52 147.655 28.52 148.655 ;
      RECT 27.52 149.655 28.52 150.655 ;
      RECT 27.52 151.655 28.52 152.655 ;
      RECT 25.52 145.655 26.52 146.655 ;
      RECT 25.52 147.655 26.52 148.655 ;
      RECT 25.52 149.655 26.52 150.655 ;
      RECT 25.52 151.655 26.52 152.655 ;
      RECT 23.52 145.655 24.52 146.655 ;
      RECT 23.52 147.655 24.52 148.655 ;
      RECT 23.52 149.655 24.52 150.655 ;
      RECT 23.52 151.655 24.52 152.655 ;
      RECT 21.52 145.655 22.52 146.655 ;
      RECT 21.52 147.655 22.52 148.655 ;
      RECT 21.52 149.655 22.52 150.655 ;
      RECT 21.52 151.655 22.52 152.655 ;
      RECT 280 142.25 290 190 ;
      RECT 240 142.25 250 190 ;
      RECT 200 60 210 190 ;
      RECT 200 142.25 290 152.25 ;
      RECT 160 43.35 170 190 ;
      RECT 70 112.9 170 122.9 ;
      RECT 70 60 80 122.9 ;
      RECT 160 43.35 203.6 53.35 ;
      RECT 90 134.45 100 190 ;
      RECT 50 134.45 60 190 ;
      RECT 10 134.45 20 190 ;
      RECT 10 134.45 100 144.45 ;
      RECT 30 60 40 144.45 ;
      RECT 215 115 225 125 ;
      RECT 209 43 219 53 ;
      RECT 21 145 29 153 ;
        RECT 10 0 20 90 ;
        RECT 50 0 60 90 ;
        RECT 90 0 100 90 ;
        RECT 220 0 230 90 ;
        RECT 0 0 350 20 ;
        RECT 140 160 150 225.2 ;
        RECT 180 160 190 207.5 ;
        RECT 140 197.5 190 207.5 ;
        RECT 260 60 270 105.55 ;
        RECT 260 95.55 330.55 105.55 ;
        RECT 320.55 95.55 330.55 219.1 ;
        RECT 0 260 350 280 ;
        RECT 240 42.165 250 90 ;
        RECT 30 160 40 250 ;
        RECT 70 160 80 250 ;
        RECT 110 160 120 250 ;
        RECT 220 160 230 250 ;
        RECT 260 160 270 208.95 ;
        RECT 300 160 310 208.95 ;
        RECT 220 198.95 310 208.95 ;
        RECT 0 230 350 250 ;
    LAYER Metal1 ;
      RECT 200 114.765 225 124.765 ;
      RECT 193.59 43.335 219 53.335 ;
      RECT 10.075 145.155 29.02 153.155 ;
  END
END MoS2Or

MACRO MoS2Xor
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MoS2Xor 0 0 ;
  SIZE 890 BY 280 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 279 27.35 291 105 ;
        RECT 19 27.35 291 39.35 ;
        RECT 239 27.35 251 95.55 ;
        RECT 39 45 51 105 ;
        RECT 19 45 51 55 ;
        RECT 19 27.35 31 205 ;
      LAYER Metal1 ;
        RECT 7.84 28.785 28.54 36.785 ;
      LAYER NSD ;
        RECT 7.84 28.785 15.84 36.785 ;
      LAYER Cont ;
        RECT 21.04 35.285 22.04 36.285 ;
        RECT 21.04 33.285 22.04 34.285 ;
        RECT 21.04 31.285 22.04 32.285 ;
        RECT 21.04 29.285 22.04 30.285 ;
        RECT 23.04 35.285 24.04 36.285 ;
        RECT 23.04 33.285 24.04 34.285 ;
        RECT 23.04 31.285 24.04 32.285 ;
        RECT 23.04 29.285 24.04 30.285 ;
        RECT 25.04 35.285 26.04 36.285 ;
        RECT 25.04 33.285 26.04 34.285 ;
        RECT 25.04 31.285 26.04 32.285 ;
        RECT 25.04 29.285 26.04 30.285 ;
        RECT 27.04 35.285 28.04 36.285 ;
        RECT 27.04 33.285 28.04 34.285 ;
        RECT 27.04 31.285 28.04 32.285 ;
        RECT 27.04 29.285 28.04 30.285 ;
      LAYER Contact ;
        RECT 8.34 35.285 9.34 36.285 ;
        RECT 8.34 33.285 9.34 34.285 ;
        RECT 8.34 31.285 9.34 32.285 ;
        RECT 8.34 29.285 9.34 30.285 ;
        RECT 10.34 35.285 11.34 36.285 ;
        RECT 10.34 33.285 11.34 34.285 ;
        RECT 10.34 31.285 11.34 32.285 ;
        RECT 10.34 29.285 11.34 30.285 ;
        RECT 12.34 35.285 13.34 36.285 ;
        RECT 12.34 33.285 13.34 34.285 ;
        RECT 12.34 31.285 13.34 32.285 ;
        RECT 12.34 29.285 13.34 30.285 ;
        RECT 14.34 35.285 15.34 36.285 ;
        RECT 14.34 33.285 15.34 34.285 ;
        RECT 14.34 31.285 15.34 32.285 ;
        RECT 14.34 29.285 15.34 30.285 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 206.6 99.25 271 111.25 ;
        RECT 259 45 271 111.25 ;
        RECT 219 45 231 111.25 ;
        RECT 39 209.65 194.65 217.65 ;
        RECT 99 45 111 105 ;
        RECT 79 45 111 55 ;
        RECT 39 122 91 134 ;
        RECT 79 45 91 134 ;
        RECT 39 122 51 217.65 ;
      LAYER Metal1 ;
        RECT 195.505 99.98 218.28 109.98 ;
        RECT 185.755 209.655 204.29 217.655 ;
        RECT 29.47 209.465 48.695 217.465 ;
      LAYER NSD ;
        RECT 195.505 99.98 205.505 217.825 ;
        RECT 29.47 209.465 37.47 217.465 ;
      LAYER Cont ;
        RECT 41.195 215.965 42.195 216.965 ;
        RECT 41.195 213.965 42.195 214.965 ;
        RECT 41.195 211.965 42.195 212.965 ;
        RECT 41.195 209.965 42.195 210.965 ;
        RECT 43.195 215.965 44.195 216.965 ;
        RECT 43.195 213.965 44.195 214.965 ;
        RECT 43.195 211.965 44.195 212.965 ;
        RECT 43.195 209.965 44.195 210.965 ;
        RECT 45.195 215.965 46.195 216.965 ;
        RECT 45.195 213.965 46.195 214.965 ;
        RECT 45.195 211.965 46.195 212.965 ;
        RECT 45.195 209.965 46.195 210.965 ;
        RECT 47.195 215.965 48.195 216.965 ;
        RECT 47.195 213.965 48.195 214.965 ;
        RECT 47.195 211.965 48.195 212.965 ;
        RECT 47.195 209.965 48.195 210.965 ;
        RECT 186.255 216.155 187.255 217.155 ;
        RECT 186.255 214.155 187.255 215.155 ;
        RECT 186.255 212.155 187.255 213.155 ;
        RECT 186.255 210.155 187.255 211.155 ;
        RECT 188.255 216.155 189.255 217.155 ;
        RECT 188.255 214.155 189.255 215.155 ;
        RECT 188.255 212.155 189.255 213.155 ;
        RECT 188.255 210.155 189.255 211.155 ;
        RECT 190.255 216.155 191.255 217.155 ;
        RECT 190.255 214.155 191.255 215.155 ;
        RECT 190.255 212.155 191.255 213.155 ;
        RECT 190.255 210.155 191.255 211.155 ;
        RECT 192.255 216.155 193.255 217.155 ;
        RECT 192.255 214.155 193.255 215.155 ;
        RECT 192.255 212.155 193.255 213.155 ;
        RECT 192.255 210.155 193.255 211.155 ;
        RECT 208.78 108.48 209.78 109.48 ;
        RECT 208.78 106.48 209.78 107.48 ;
        RECT 208.78 104.48 209.78 105.48 ;
        RECT 208.78 102.48 209.78 103.48 ;
        RECT 208.78 100.48 209.78 101.48 ;
        RECT 210.78 108.48 211.78 109.48 ;
        RECT 210.78 106.48 211.78 107.48 ;
        RECT 210.78 104.48 211.78 105.48 ;
        RECT 210.78 102.48 211.78 103.48 ;
        RECT 210.78 100.48 211.78 101.48 ;
        RECT 212.78 108.48 213.78 109.48 ;
        RECT 212.78 106.48 213.78 107.48 ;
        RECT 212.78 104.48 213.78 105.48 ;
        RECT 212.78 102.48 213.78 103.48 ;
        RECT 212.78 100.48 213.78 101.48 ;
        RECT 214.78 108.48 215.78 109.48 ;
        RECT 214.78 106.48 215.78 107.48 ;
        RECT 214.78 104.48 215.78 105.48 ;
        RECT 214.78 102.48 215.78 103.48 ;
        RECT 214.78 100.48 215.78 101.48 ;
        RECT 216.78 108.48 217.78 109.48 ;
        RECT 216.78 106.48 217.78 107.48 ;
        RECT 216.78 104.48 217.78 105.48 ;
        RECT 216.78 102.48 217.78 103.48 ;
        RECT 216.78 100.48 217.78 101.48 ;
      LAYER Contact ;
        RECT 29.97 215.965 30.97 216.965 ;
        RECT 29.97 213.965 30.97 214.965 ;
        RECT 29.97 211.965 30.97 212.965 ;
        RECT 29.97 209.965 30.97 210.965 ;
        RECT 31.97 215.965 32.97 216.965 ;
        RECT 31.97 213.965 32.97 214.965 ;
        RECT 31.97 211.965 32.97 212.965 ;
        RECT 31.97 209.965 32.97 210.965 ;
        RECT 33.97 215.965 34.97 216.965 ;
        RECT 33.97 213.965 34.97 214.965 ;
        RECT 33.97 211.965 34.97 212.965 ;
        RECT 33.97 209.965 34.97 210.965 ;
        RECT 35.97 215.965 36.97 216.965 ;
        RECT 35.97 213.965 36.97 214.965 ;
        RECT 35.97 211.965 36.97 212.965 ;
        RECT 35.97 209.965 36.97 210.965 ;
        RECT 196.005 108.48 197.005 109.48 ;
        RECT 196.005 106.48 197.005 107.48 ;
        RECT 196.005 104.48 197.005 105.48 ;
        RECT 196.005 102.48 197.005 103.48 ;
        RECT 196.005 100.48 197.005 101.48 ;
        RECT 196.79 216.155 197.79 217.155 ;
        RECT 196.79 214.155 197.79 215.155 ;
        RECT 196.79 212.155 197.79 213.155 ;
        RECT 196.79 210.155 197.79 211.155 ;
        RECT 198.005 108.48 199.005 109.48 ;
        RECT 198.005 106.48 199.005 107.48 ;
        RECT 198.005 104.48 199.005 105.48 ;
        RECT 198.005 102.48 199.005 103.48 ;
        RECT 198.005 100.48 199.005 101.48 ;
        RECT 198.79 216.155 199.79 217.155 ;
        RECT 198.79 214.155 199.79 215.155 ;
        RECT 198.79 212.155 199.79 213.155 ;
        RECT 198.79 210.155 199.79 211.155 ;
        RECT 200.005 108.48 201.005 109.48 ;
        RECT 200.005 106.48 201.005 107.48 ;
        RECT 200.005 104.48 201.005 105.48 ;
        RECT 200.005 102.48 201.005 103.48 ;
        RECT 200.005 100.48 201.005 101.48 ;
        RECT 200.79 216.155 201.79 217.155 ;
        RECT 200.79 214.155 201.79 215.155 ;
        RECT 200.79 212.155 201.79 213.155 ;
        RECT 200.79 210.155 201.79 211.155 ;
        RECT 202.005 108.48 203.005 109.48 ;
        RECT 202.005 106.48 203.005 107.48 ;
        RECT 202.005 104.48 203.005 105.48 ;
        RECT 202.005 102.48 203.005 103.48 ;
        RECT 202.005 100.48 203.005 101.48 ;
        RECT 202.79 216.155 203.79 217.155 ;
        RECT 202.79 214.155 203.79 215.155 ;
        RECT 202.79 212.155 203.79 213.155 ;
        RECT 202.79 210.155 203.79 211.155 ;
        RECT 204.005 108.48 205.005 109.48 ;
        RECT 204.005 106.48 205.005 107.48 ;
        RECT 204.005 104.48 205.005 105.48 ;
        RECT 204.005 102.48 205.005 103.48 ;
        RECT 204.005 100.48 205.005 101.48 ;
    END
  END B
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 10 42.95 20 190 ;
    END
    PORT
      LAYER NSD ;
        RECT 10 42.95 60 52.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 50 0 60 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 210 0 220 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 250 0 260 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 290 0 300 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 420 0 430 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 560 0 570 190 ;
    END
    PORT
      LAYER NSD ;
        RECT 600 0 610 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 750 0 760 90 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 0 890 20 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Contact ;
        RECT 863 211.225 864 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 863 213.225 864 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 863 215.225 864 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 863 217.225 864 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 863 261.65 864 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 863 263.65 864 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 863 265.65 864 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 863 267.65 864 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 861 211.225 862 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 861 213.225 862 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 861 215.225 862 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 861 217.225 862 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 861 261.65 862 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 861 263.65 862 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 861 265.65 862 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 861 267.65 862 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 859 211.225 860 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 859 213.225 860 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 859 215.225 860 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 859 217.225 860 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 859 261.65 860 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 859 263.65 860 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 859 265.65 860 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 859 267.65 860 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 857 211.225 858 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 857 213.225 858 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 857 215.225 858 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 857 217.225 858 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 857 261.65 858 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 857 263.65 858 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 857 265.65 858 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 857 267.65 858 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 721.465 212.915 722.465 213.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 721.465 214.915 722.465 215.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 721.465 216.915 722.465 217.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 721.465 218.915 722.465 219.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 721.465 261.91 722.465 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 721.465 263.91 722.465 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 721.465 265.91 722.465 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 721.465 267.91 722.465 268.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 719.465 212.915 720.465 213.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 719.465 214.915 720.465 215.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 719.465 216.915 720.465 217.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 719.465 218.915 720.465 219.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 719.465 261.91 720.465 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 719.465 263.91 720.465 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 719.465 265.91 720.465 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 719.465 267.91 720.465 268.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 717.465 212.915 718.465 213.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 717.465 214.915 718.465 215.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 717.465 216.915 718.465 217.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 717.465 218.915 718.465 219.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 717.465 261.91 718.465 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 717.465 263.91 718.465 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 717.465 265.91 718.465 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 717.465 267.91 718.465 268.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 715.465 212.915 716.465 213.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 715.465 214.915 716.465 215.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 715.465 216.915 716.465 217.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 715.465 218.915 716.465 219.915 ;
    END
    PORT
      LAYER Contact ;
        RECT 715.465 261.91 716.465 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 715.465 263.91 716.465 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 715.465 265.91 716.465 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 715.465 267.91 716.465 268.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 528.2 211.225 529.2 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 528.2 213.225 529.2 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 528.2 215.225 529.2 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 528.2 217.225 529.2 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 528.2 261.65 529.2 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 528.2 263.65 529.2 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 528.2 265.65 529.2 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 528.2 267.65 529.2 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 526.2 211.225 527.2 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 526.2 213.225 527.2 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 526.2 215.225 527.2 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 526.2 217.225 527.2 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 526.2 261.65 527.2 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 526.2 263.65 527.2 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 526.2 265.65 527.2 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 526.2 267.65 527.2 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 524.2 211.225 525.2 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 524.2 213.225 525.2 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 524.2 215.225 525.2 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 524.2 217.225 525.2 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 524.2 261.65 525.2 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 524.2 263.65 525.2 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 524.2 265.65 525.2 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 524.2 267.65 525.2 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 522.2 211.225 523.2 212.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 522.2 213.225 523.2 214.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 522.2 215.225 523.2 216.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 522.2 217.225 523.2 218.225 ;
    END
    PORT
      LAYER Contact ;
        RECT 522.2 261.65 523.2 262.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 522.2 263.65 523.2 264.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 522.2 265.65 523.2 266.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 522.2 267.65 523.2 268.65 ;
    END
    PORT
      LAYER Contact ;
        RECT 347.445 216.875 348.445 217.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 347.445 218.875 348.445 219.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 347.445 220.875 348.445 221.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 347.445 222.875 348.445 223.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 347.445 262.575 348.445 263.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 347.445 264.575 348.445 265.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 347.445 266.575 348.445 267.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 347.445 268.575 348.445 269.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 345.445 216.875 346.445 217.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 345.445 218.875 346.445 219.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 345.445 220.875 346.445 221.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 345.445 222.875 346.445 223.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 345.445 262.575 346.445 263.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 345.445 264.575 346.445 265.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 345.445 266.575 346.445 267.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 345.445 268.575 346.445 269.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 343.445 216.875 344.445 217.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 343.445 218.875 344.445 219.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 343.445 220.875 344.445 221.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 343.445 222.875 344.445 223.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 343.445 262.575 344.445 263.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 343.445 264.575 344.445 265.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 343.445 266.575 344.445 267.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 343.445 268.575 344.445 269.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 341.445 216.875 342.445 217.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 341.445 218.875 342.445 219.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 341.445 220.875 342.445 221.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 341.445 222.875 342.445 223.875 ;
    END
    PORT
      LAYER Contact ;
        RECT 341.445 262.575 342.445 263.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 341.445 264.575 342.445 265.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 341.445 266.575 342.445 267.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 341.445 268.575 342.445 269.575 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.26 219.77 174.26 220.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.26 221.77 174.26 222.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.26 223.77 174.26 224.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.26 225.77 174.26 226.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.26 261.91 174.26 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.26 263.91 174.26 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.26 265.91 174.26 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 173.26 267.91 174.26 268.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.26 219.77 172.26 220.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.26 221.77 172.26 222.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.26 223.77 172.26 224.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.26 225.77 172.26 226.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.26 261.91 172.26 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.26 263.91 172.26 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.26 265.91 172.26 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 171.26 267.91 172.26 268.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.26 219.77 170.26 220.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.26 221.77 170.26 222.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.26 223.77 170.26 224.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.26 225.77 170.26 226.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.26 261.91 170.26 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.26 263.91 170.26 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.26 265.91 170.26 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 169.26 267.91 170.26 268.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.26 219.77 168.26 220.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.26 221.77 168.26 222.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.26 223.77 168.26 224.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.26 225.77 168.26 226.77 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.26 261.91 168.26 262.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.26 263.91 168.26 264.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.26 265.91 168.26 266.91 ;
    END
    PORT
      LAYER Contact ;
        RECT 167.26 267.91 168.26 268.91 ;
    END
    PORT
      LAYER NSD ;
        RECT 150 60 160 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 150 98.9 175.7 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 165.7 98.9 175.7 227.35 ;
    END
    PORT
      LAYER NSD ;
        RECT 340 160 350 225.2 ;
    END
    PORT
      LAYER NSD ;
        RECT 380 160 390 207.5 ;
    END
    PORT
      LAYER NSD ;
        RECT 340 197.5 390 207.5 ;
    END
    PORT
      LAYER NSD ;
        RECT 460 60 470 105.55 ;
    END
    PORT
      LAYER NSD ;
        RECT 460 95.55 530.55 105.55 ;
    END
    PORT
      LAYER NSD ;
        RECT 520.55 95.55 530.55 219.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 700 60 710 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 700 98.9 723.85 108.9 ;
    END
    PORT
      LAYER NSD ;
        RECT 713.85 98.9 723.85 220.75 ;
    END
    PORT
      LAYER NSD ;
        RECT 790 60 800 105.55 ;
    END
    PORT
      LAYER NSD ;
        RECT 790 95.55 865.45 105.55 ;
    END
    PORT
      LAYER NSD ;
        RECT 855.45 95.55 865.45 219.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 260 890 280 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 166.76 219.27 174.76 269.41 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 340.945 216.375 348.945 270.075 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 521.7 210.725 529.7 269.15 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 714.965 212.415 722.965 269.41 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 856.5 210.725 864.5 269.15 ;
    END
  END VDD
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER NSD ;
        RECT 770 31.785 780 90 ;
    END
  END VOUT
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 70 160 80 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 110 160 120 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 150 160 160 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 70 198.1 160 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 230 160 240 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 270 160 280 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 310 160 320 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 420 160 430 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 460 160 470 208.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 500 160 510 208.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 420 198.95 510 208.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 620 160 630 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 660 160 670 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 700 160 710 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 620 198.1 710 208.1 ;
    END
    PORT
      LAYER NSD ;
        RECT 750 160 760 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 790 160 800 208.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 830 160 840 208.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 750 198.95 840 208.95 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 230 890 250 ;
    END
  END VSS
  OBS
    LAYER Gate ;
      RECT 799 195 831 205 ;
      RECT 819 145 831 205 ;
      RECT 759 195 791 205 ;
      RECT 779 45 791 205 ;
      RECT 739 145 751 205 ;
      RECT 799 145 811 205 ;
      RECT 759 145 771 205 ;
      RECT 779 145 811 155 ;
      RECT 739 145 771 155 ;
      RECT 745 114.75 791 124.75 ;
      RECT 759 43.35 771 105 ;
      RECT 739 43.35 751 105 ;
      RECT 739 43.35 771 55.35 ;
      RECT 669 195 701 205 ;
      RECT 689 145 701 205 ;
      RECT 629 195 661 205 ;
      RECT 649 145 661 205 ;
      RECT 609 145 621 205 ;
      RECT 669 122.6 681 205 ;
      RECT 629 145 641 205 ;
      RECT 649 145 681 155 ;
      RECT 609 145 641 155 ;
      RECT 669 122.6 701 134.6 ;
      RECT 689 45 701 134.6 ;
      RECT 534.6 210.1 601 222.1 ;
      RECT 589 122 601 222.1 ;
      RECT 589 122 641 134 ;
      RECT 629 45 641 134 ;
      RECT 649 45 661 105 ;
      RECT 629 45 661 55 ;
      RECT 569 21.45 581 205 ;
      RECT 589 45 601 105 ;
      RECT 569 45 601 55 ;
      RECT 440.1 21.45 581 33.45 ;
      RECT 469 195 501 205 ;
      RECT 489 145 501 205 ;
      RECT 429 195 461 205 ;
      RECT 449 45 461 205 ;
      RECT 409 145 421 205 ;
      RECT 469 145 481 205 ;
      RECT 429 145 441 205 ;
      RECT 449 145 481 155 ;
      RECT 409 145 441 155 ;
      RECT 415 114.75 461 124.75 ;
      RECT 429 44.95 441 105 ;
      RECT 409 44.95 421 105 ;
      RECT 373.55 44.95 441 56.95 ;
      RECT 369 145 381 205 ;
      RECT 279 195 361 205 ;
      RECT 349 145 361 205 ;
      RECT 239 195 271 205 ;
      RECT 259 145 271 205 ;
      RECT 219 145 231 205 ;
      RECT 299 193 361 205 ;
      RECT 279 145 291 205 ;
      RECT 239 145 251 205 ;
      RECT 299 145 311 205 ;
      RECT 349 145 381 155 ;
      RECT 259 145 291 155 ;
      RECT 219 145 251 155 ;
      RECT 119 195 151 205 ;
      RECT 139 145 151 205 ;
      RECT 79 195 111 205 ;
      RECT 99 145 111 205 ;
      RECT 59 145 71 205 ;
      RECT 119 122.6 131 205 ;
      RECT 79 145 91 205 ;
      RECT 99 145 131 155 ;
      RECT 59 145 91 155 ;
      RECT 119 122.6 151 134.6 ;
      RECT 139 45 151 134.6 ;
    LAYER NSD ;
      RECT 810 142.25 820 190 ;
      RECT 770 142.25 780 190 ;
      RECT 730 60 740 190 ;
      RECT 730 142.25 820 152.25 ;
      RECT 640 96.35 690 106.35 ;
      RECT 680 43.35 690 106.35 ;
      RECT 640 60 650 106.35 ;
      RECT 680 43.35 733.15 53.35 ;
      RECT 680 141.75 690 190 ;
      RECT 640 141.75 650 190 ;
      RECT 600 141.75 610 190 ;
      RECT 600 141.75 690 151.75 ;
      RECT 658.6 131.2 666.6 151.75 ;
      RECT 580 96.35 630 106.35 ;
      RECT 620 42.05 630 106.35 ;
      RECT 580 60 590 106.35 ;
      RECT 660 42.05 670 90 ;
      RECT 620 42.05 670 52.05 ;
      RECT 480 142.25 490 190 ;
      RECT 440 142.25 450 190 ;
      RECT 400 60 410 190 ;
      RECT 400 142.25 490 152.25 ;
      RECT 360 45.85 370 190 ;
      RECT 270 112.9 370 122.9 ;
      RECT 270 60 280 122.9 ;
      RECT 290 134.45 300 190 ;
      RECT 250 134.45 260 190 ;
      RECT 210 134.45 220 190 ;
      RECT 210 134.45 300 144.45 ;
      RECT 230 60 240 144.45 ;
      RECT 90 96.35 140 106.35 ;
      RECT 130 43.4 140 106.35 ;
      RECT 90 60 100 106.35 ;
      RECT 130 141.75 140 190 ;
      RECT 90 141.75 100 190 ;
      RECT 50 141.75 60 190 ;
      RECT 50 141.75 140 151.75 ;
      RECT 108.6 131.2 116.6 151.75 ;
      RECT 30 96.35 80 106.35 ;
      RECT 70 42.05 80 106.35 ;
      RECT 30 60 40 106.35 ;
      RECT 110 42.05 120 90 ;
      RECT 70 42.05 120 52.05 ;
      RECT 580 160 590 190 ;
      RECT 536.575 46.185 544.575 207.105 ;
      RECT 440 34.505 450 90 ;
      RECT 30 160 40 190 ;
    LAYER Contact ;
      RECT 738.5 115.265 739.5 116.265 ;
      RECT 738.5 117.265 739.5 118.265 ;
      RECT 738.5 119.265 739.5 120.265 ;
      RECT 738.5 121.265 739.5 122.265 ;
      RECT 738.5 123.265 739.5 124.265 ;
      RECT 736.5 115.265 737.5 116.265 ;
      RECT 736.5 117.265 737.5 118.265 ;
      RECT 736.5 119.265 737.5 120.265 ;
      RECT 736.5 121.265 737.5 122.265 ;
      RECT 736.5 123.265 737.5 124.265 ;
      RECT 734.5 115.265 735.5 116.265 ;
      RECT 734.5 117.265 735.5 118.265 ;
      RECT 734.5 119.265 735.5 120.265 ;
      RECT 734.5 121.265 735.5 122.265 ;
      RECT 734.5 123.265 735.5 124.265 ;
      RECT 732.5 115.265 733.5 116.265 ;
      RECT 732.5 117.265 733.5 118.265 ;
      RECT 732.5 119.265 733.5 120.265 ;
      RECT 732.5 121.265 733.5 122.265 ;
      RECT 732.5 123.265 733.5 124.265 ;
      RECT 731.665 43.835 732.665 44.835 ;
      RECT 731.665 45.835 732.665 46.835 ;
      RECT 731.665 47.835 732.665 48.835 ;
      RECT 731.665 49.835 732.665 50.835 ;
      RECT 731.665 51.835 732.665 52.835 ;
      RECT 730.5 115.265 731.5 116.265 ;
      RECT 730.5 117.265 731.5 118.265 ;
      RECT 730.5 119.265 731.5 120.265 ;
      RECT 730.5 121.265 731.5 122.265 ;
      RECT 730.5 123.265 731.5 124.265 ;
      RECT 729.665 43.835 730.665 44.835 ;
      RECT 729.665 45.835 730.665 46.835 ;
      RECT 729.665 47.835 730.665 48.835 ;
      RECT 729.665 49.835 730.665 50.835 ;
      RECT 729.665 51.835 730.665 52.835 ;
      RECT 727.665 43.835 728.665 44.835 ;
      RECT 727.665 45.835 728.665 46.835 ;
      RECT 727.665 47.835 728.665 48.835 ;
      RECT 727.665 49.835 728.665 50.835 ;
      RECT 727.665 51.835 728.665 52.835 ;
      RECT 725.665 43.835 726.665 44.835 ;
      RECT 725.665 45.835 726.665 46.835 ;
      RECT 725.665 47.835 726.665 48.835 ;
      RECT 725.665 49.835 726.665 50.835 ;
      RECT 725.665 51.835 726.665 52.835 ;
      RECT 723.665 43.835 724.665 44.835 ;
      RECT 723.665 45.835 724.665 46.835 ;
      RECT 723.665 47.835 724.665 48.835 ;
      RECT 723.665 49.835 724.665 50.835 ;
      RECT 723.665 51.835 724.665 52.835 ;
      RECT 665.11 131.675 666.11 132.675 ;
      RECT 665.11 133.675 666.11 134.675 ;
      RECT 665.11 135.675 666.11 136.675 ;
      RECT 665.11 137.675 666.11 138.675 ;
      RECT 663.11 131.675 664.11 132.675 ;
      RECT 663.11 133.675 664.11 134.675 ;
      RECT 663.11 135.675 664.11 136.675 ;
      RECT 663.11 137.675 664.11 138.675 ;
      RECT 661.11 131.675 662.11 132.675 ;
      RECT 661.11 133.675 662.11 134.675 ;
      RECT 661.11 135.675 662.11 136.675 ;
      RECT 661.11 137.675 662.11 138.675 ;
      RECT 659.11 131.675 660.11 132.675 ;
      RECT 659.11 133.675 660.11 134.675 ;
      RECT 659.11 135.675 660.11 136.675 ;
      RECT 659.11 137.675 660.11 138.675 ;
      RECT 543.075 46.685 544.075 47.685 ;
      RECT 543.075 48.685 544.075 49.685 ;
      RECT 543.075 50.685 544.075 51.685 ;
      RECT 543.075 52.685 544.075 53.685 ;
      RECT 543.075 199.605 544.075 200.605 ;
      RECT 543.075 201.605 544.075 202.605 ;
      RECT 543.075 203.605 544.075 204.605 ;
      RECT 543.075 205.605 544.075 206.605 ;
      RECT 541.075 46.685 542.075 47.685 ;
      RECT 541.075 48.685 542.075 49.685 ;
      RECT 541.075 50.685 542.075 51.685 ;
      RECT 541.075 52.685 542.075 53.685 ;
      RECT 541.075 199.605 542.075 200.605 ;
      RECT 541.075 201.605 542.075 202.605 ;
      RECT 541.075 203.605 542.075 204.605 ;
      RECT 541.075 205.605 542.075 206.605 ;
      RECT 539.075 46.685 540.075 47.685 ;
      RECT 539.075 48.685 540.075 49.685 ;
      RECT 539.075 50.685 540.075 51.685 ;
      RECT 539.075 52.685 540.075 53.685 ;
      RECT 539.075 199.605 540.075 200.605 ;
      RECT 539.075 201.605 540.075 202.605 ;
      RECT 539.075 203.605 540.075 204.605 ;
      RECT 539.075 205.605 540.075 206.605 ;
      RECT 537.075 46.685 538.075 47.685 ;
      RECT 537.075 48.685 538.075 49.685 ;
      RECT 537.075 50.685 538.075 51.685 ;
      RECT 537.075 52.685 538.075 53.685 ;
      RECT 537.075 199.605 538.075 200.605 ;
      RECT 537.075 201.605 538.075 202.605 ;
      RECT 537.075 203.605 538.075 204.605 ;
      RECT 537.075 205.605 538.075 206.605 ;
      RECT 447.785 36.005 448.785 37.005 ;
      RECT 447.785 38.005 448.785 39.005 ;
      RECT 447.785 40.005 448.785 41.005 ;
      RECT 447.785 42.005 448.785 43.005 ;
      RECT 445.785 36.005 446.785 37.005 ;
      RECT 445.785 38.005 446.785 39.005 ;
      RECT 445.785 40.005 446.785 41.005 ;
      RECT 445.785 42.005 446.785 43.005 ;
      RECT 443.785 36.005 444.785 37.005 ;
      RECT 443.785 38.005 444.785 39.005 ;
      RECT 443.785 40.005 444.785 41.005 ;
      RECT 443.785 42.005 444.785 43.005 ;
      RECT 441.785 36.005 442.785 37.005 ;
      RECT 441.785 38.005 442.785 39.005 ;
      RECT 441.785 40.005 442.785 41.005 ;
      RECT 441.785 42.005 442.785 43.005 ;
      RECT 408.5 115.265 409.5 116.265 ;
      RECT 408.5 117.265 409.5 118.265 ;
      RECT 408.5 119.265 409.5 120.265 ;
      RECT 408.5 121.265 409.5 122.265 ;
      RECT 408.5 123.265 409.5 124.265 ;
      RECT 406.5 115.265 407.5 116.265 ;
      RECT 406.5 117.265 407.5 118.265 ;
      RECT 406.5 119.265 407.5 120.265 ;
      RECT 406.5 121.265 407.5 122.265 ;
      RECT 406.5 123.265 407.5 124.265 ;
      RECT 404.5 115.265 405.5 116.265 ;
      RECT 404.5 117.265 405.5 118.265 ;
      RECT 404.5 119.265 405.5 120.265 ;
      RECT 404.5 121.265 405.5 122.265 ;
      RECT 404.5 123.265 405.5 124.265 ;
      RECT 402.5 115.265 403.5 116.265 ;
      RECT 402.5 117.265 403.5 118.265 ;
      RECT 402.5 119.265 403.5 120.265 ;
      RECT 402.5 121.265 403.5 122.265 ;
      RECT 402.5 123.265 403.5 124.265 ;
      RECT 400.5 115.265 401.5 116.265 ;
      RECT 400.5 117.265 401.5 118.265 ;
      RECT 400.5 119.265 401.5 120.265 ;
      RECT 400.5 121.265 401.5 122.265 ;
      RECT 400.5 123.265 401.5 124.265 ;
      RECT 368.5 46.76 369.5 47.76 ;
      RECT 368.5 48.76 369.5 49.76 ;
      RECT 368.5 50.76 369.5 51.76 ;
      RECT 368.5 52.76 369.5 53.76 ;
      RECT 368.5 54.76 369.5 55.76 ;
      RECT 366.5 46.76 367.5 47.76 ;
      RECT 366.5 48.76 367.5 49.76 ;
      RECT 366.5 50.76 367.5 51.76 ;
      RECT 366.5 52.76 367.5 53.76 ;
      RECT 366.5 54.76 367.5 55.76 ;
      RECT 364.5 46.76 365.5 47.76 ;
      RECT 364.5 48.76 365.5 49.76 ;
      RECT 364.5 50.76 365.5 51.76 ;
      RECT 364.5 52.76 365.5 53.76 ;
      RECT 364.5 54.76 365.5 55.76 ;
      RECT 362.5 46.76 363.5 47.76 ;
      RECT 362.5 48.76 363.5 49.76 ;
      RECT 362.5 50.76 363.5 51.76 ;
      RECT 362.5 52.76 363.5 53.76 ;
      RECT 362.5 54.76 363.5 55.76 ;
      RECT 360.5 46.76 361.5 47.76 ;
      RECT 360.5 48.76 361.5 49.76 ;
      RECT 360.5 50.76 361.5 51.76 ;
      RECT 360.5 52.76 361.5 53.76 ;
      RECT 360.5 54.76 361.5 55.76 ;
      RECT 216.575 145.655 217.575 146.655 ;
      RECT 216.575 147.655 217.575 148.655 ;
      RECT 216.575 149.655 217.575 150.655 ;
      RECT 216.575 151.655 217.575 152.655 ;
      RECT 214.575 145.655 215.575 146.655 ;
      RECT 214.575 147.655 215.575 148.655 ;
      RECT 214.575 149.655 215.575 150.655 ;
      RECT 214.575 151.655 215.575 152.655 ;
      RECT 212.575 145.655 213.575 146.655 ;
      RECT 212.575 147.655 213.575 148.655 ;
      RECT 212.575 149.655 213.575 150.655 ;
      RECT 212.575 151.655 213.575 152.655 ;
      RECT 210.575 145.655 211.575 146.655 ;
      RECT 210.575 147.655 211.575 148.655 ;
      RECT 210.575 149.655 211.575 150.655 ;
      RECT 210.575 151.655 211.575 152.655 ;
      RECT 136.78 44.125 137.78 45.125 ;
      RECT 136.78 46.125 137.78 47.125 ;
      RECT 136.78 48.125 137.78 49.125 ;
      RECT 136.78 50.125 137.78 51.125 ;
      RECT 134.78 44.125 135.78 45.125 ;
      RECT 134.78 46.125 135.78 47.125 ;
      RECT 134.78 48.125 135.78 49.125 ;
      RECT 134.78 50.125 135.78 51.125 ;
      RECT 132.78 44.125 133.78 45.125 ;
      RECT 132.78 46.125 133.78 47.125 ;
      RECT 132.78 48.125 133.78 49.125 ;
      RECT 132.78 50.125 133.78 51.125 ;
      RECT 130.78 44.125 131.78 45.125 ;
      RECT 130.78 46.125 131.78 47.125 ;
      RECT 130.78 48.125 131.78 49.125 ;
      RECT 130.78 50.125 131.78 51.125 ;
      RECT 115.11 131.675 116.11 132.675 ;
      RECT 115.11 133.675 116.11 134.675 ;
      RECT 115.11 135.675 116.11 136.675 ;
      RECT 115.11 137.675 116.11 138.675 ;
      RECT 113.11 131.675 114.11 132.675 ;
      RECT 113.11 133.675 114.11 134.675 ;
      RECT 113.11 135.675 114.11 136.675 ;
      RECT 113.11 137.675 114.11 138.675 ;
      RECT 111.11 131.675 112.11 132.675 ;
      RECT 111.11 133.675 112.11 134.675 ;
      RECT 111.11 135.675 112.11 136.675 ;
      RECT 111.11 137.675 112.11 138.675 ;
      RECT 109.11 131.675 110.11 132.675 ;
      RECT 109.11 133.675 110.11 134.675 ;
      RECT 109.11 135.675 110.11 136.675 ;
      RECT 109.11 137.675 110.11 138.675 ;
    LAYER Cont ;
      RECT 753.5 115.265 754.5 116.265 ;
      RECT 753.5 117.265 754.5 118.265 ;
      RECT 753.5 119.265 754.5 120.265 ;
      RECT 753.5 121.265 754.5 122.265 ;
      RECT 753.5 123.265 754.5 124.265 ;
      RECT 751.5 115.265 752.5 116.265 ;
      RECT 751.5 117.265 752.5 118.265 ;
      RECT 751.5 119.265 752.5 120.265 ;
      RECT 751.5 121.265 752.5 122.265 ;
      RECT 751.5 123.265 752.5 124.265 ;
      RECT 749.5 115.265 750.5 116.265 ;
      RECT 749.5 117.265 750.5 118.265 ;
      RECT 749.5 119.265 750.5 120.265 ;
      RECT 749.5 121.265 750.5 122.265 ;
      RECT 749.5 123.265 750.5 124.265 ;
      RECT 747.5 43.835 748.5 44.835 ;
      RECT 747.5 45.835 748.5 46.835 ;
      RECT 747.5 47.835 748.5 48.835 ;
      RECT 747.5 49.835 748.5 50.835 ;
      RECT 747.5 51.835 748.5 52.835 ;
      RECT 747.5 115.265 748.5 116.265 ;
      RECT 747.5 117.265 748.5 118.265 ;
      RECT 747.5 119.265 748.5 120.265 ;
      RECT 747.5 121.265 748.5 122.265 ;
      RECT 747.5 123.265 748.5 124.265 ;
      RECT 745.5 43.835 746.5 44.835 ;
      RECT 745.5 45.835 746.5 46.835 ;
      RECT 745.5 47.835 746.5 48.835 ;
      RECT 745.5 49.835 746.5 50.835 ;
      RECT 745.5 51.835 746.5 52.835 ;
      RECT 745.5 115.265 746.5 116.265 ;
      RECT 745.5 117.265 746.5 118.265 ;
      RECT 745.5 119.265 746.5 120.265 ;
      RECT 745.5 121.265 746.5 122.265 ;
      RECT 745.5 123.265 746.5 124.265 ;
      RECT 743.5 43.835 744.5 44.835 ;
      RECT 743.5 45.835 744.5 46.835 ;
      RECT 743.5 47.835 744.5 48.835 ;
      RECT 743.5 49.835 744.5 50.835 ;
      RECT 743.5 51.835 744.5 52.835 ;
      RECT 741.5 43.835 742.5 44.835 ;
      RECT 741.5 45.835 742.5 46.835 ;
      RECT 741.5 47.835 742.5 48.835 ;
      RECT 741.5 49.835 742.5 50.835 ;
      RECT 741.5 51.835 742.5 52.835 ;
      RECT 739.5 43.835 740.5 44.835 ;
      RECT 739.5 45.835 740.5 46.835 ;
      RECT 739.5 47.835 740.5 48.835 ;
      RECT 739.5 49.835 740.5 50.835 ;
      RECT 739.5 51.835 740.5 52.835 ;
      RECT 676.925 131.675 677.925 132.675 ;
      RECT 676.925 133.675 677.925 134.675 ;
      RECT 676.925 135.675 677.925 136.675 ;
      RECT 676.925 137.675 677.925 138.675 ;
      RECT 674.925 131.675 675.925 132.675 ;
      RECT 674.925 133.675 675.925 134.675 ;
      RECT 674.925 135.675 675.925 136.675 ;
      RECT 674.925 137.675 675.925 138.675 ;
      RECT 672.925 131.675 673.925 132.675 ;
      RECT 672.925 133.675 673.925 134.675 ;
      RECT 672.925 135.675 673.925 136.675 ;
      RECT 672.925 137.675 673.925 138.675 ;
      RECT 670.925 131.675 671.925 132.675 ;
      RECT 670.925 133.675 671.925 134.675 ;
      RECT 670.925 135.675 671.925 136.675 ;
      RECT 670.925 137.675 671.925 138.675 ;
      RECT 543.075 210.83 544.075 211.83 ;
      RECT 543.075 212.83 544.075 213.83 ;
      RECT 543.075 214.83 544.075 215.83 ;
      RECT 543.075 216.83 544.075 217.83 ;
      RECT 541.075 210.83 542.075 211.83 ;
      RECT 541.075 212.83 542.075 213.83 ;
      RECT 541.075 214.83 542.075 215.83 ;
      RECT 541.075 216.83 542.075 217.83 ;
      RECT 539.075 210.83 540.075 211.83 ;
      RECT 539.075 212.83 540.075 213.83 ;
      RECT 539.075 214.83 540.075 215.83 ;
      RECT 539.075 216.83 540.075 217.83 ;
      RECT 537.075 210.83 538.075 211.83 ;
      RECT 537.075 212.83 538.075 213.83 ;
      RECT 537.075 214.83 538.075 215.83 ;
      RECT 537.075 216.83 538.075 217.83 ;
      RECT 447.785 23.305 448.785 24.305 ;
      RECT 447.785 25.305 448.785 26.305 ;
      RECT 447.785 27.305 448.785 28.305 ;
      RECT 447.785 29.305 448.785 30.305 ;
      RECT 445.785 23.305 446.785 24.305 ;
      RECT 445.785 25.305 446.785 26.305 ;
      RECT 445.785 27.305 446.785 28.305 ;
      RECT 445.785 29.305 446.785 30.305 ;
      RECT 443.785 23.305 444.785 24.305 ;
      RECT 443.785 25.305 444.785 26.305 ;
      RECT 443.785 27.305 444.785 28.305 ;
      RECT 443.785 29.305 444.785 30.305 ;
      RECT 441.785 23.305 442.785 24.305 ;
      RECT 441.785 25.305 442.785 26.305 ;
      RECT 441.785 27.305 442.785 28.305 ;
      RECT 441.785 29.305 442.785 30.305 ;
      RECT 423.5 115.265 424.5 116.265 ;
      RECT 423.5 117.265 424.5 118.265 ;
      RECT 423.5 119.265 424.5 120.265 ;
      RECT 423.5 121.265 424.5 122.265 ;
      RECT 423.5 123.265 424.5 124.265 ;
      RECT 421.5 115.265 422.5 116.265 ;
      RECT 421.5 117.265 422.5 118.265 ;
      RECT 421.5 119.265 422.5 120.265 ;
      RECT 421.5 121.265 422.5 122.265 ;
      RECT 421.5 123.265 422.5 124.265 ;
      RECT 419.5 115.265 420.5 116.265 ;
      RECT 419.5 117.265 420.5 118.265 ;
      RECT 419.5 119.265 420.5 120.265 ;
      RECT 419.5 121.265 420.5 122.265 ;
      RECT 419.5 123.265 420.5 124.265 ;
      RECT 417.5 115.265 418.5 116.265 ;
      RECT 417.5 117.265 418.5 118.265 ;
      RECT 417.5 119.265 418.5 120.265 ;
      RECT 417.5 121.265 418.5 122.265 ;
      RECT 417.5 123.265 418.5 124.265 ;
      RECT 415.5 115.265 416.5 116.265 ;
      RECT 415.5 117.265 416.5 118.265 ;
      RECT 415.5 119.265 416.5 120.265 ;
      RECT 415.5 121.265 416.5 122.265 ;
      RECT 415.5 123.265 416.5 124.265 ;
      RECT 382.525 46.76 383.525 47.76 ;
      RECT 382.525 48.76 383.525 49.76 ;
      RECT 382.525 50.76 383.525 51.76 ;
      RECT 382.525 52.76 383.525 53.76 ;
      RECT 382.525 54.76 383.525 55.76 ;
      RECT 380.525 46.76 381.525 47.76 ;
      RECT 380.525 48.76 381.525 49.76 ;
      RECT 380.525 50.76 381.525 51.76 ;
      RECT 380.525 52.76 381.525 53.76 ;
      RECT 380.525 54.76 381.525 55.76 ;
      RECT 378.525 46.76 379.525 47.76 ;
      RECT 378.525 48.76 379.525 49.76 ;
      RECT 378.525 50.76 379.525 51.76 ;
      RECT 378.525 52.76 379.525 53.76 ;
      RECT 378.525 54.76 379.525 55.76 ;
      RECT 376.525 46.76 377.525 47.76 ;
      RECT 376.525 48.76 377.525 49.76 ;
      RECT 376.525 50.76 377.525 51.76 ;
      RECT 376.525 52.76 377.525 53.76 ;
      RECT 376.525 54.76 377.525 55.76 ;
      RECT 374.525 46.76 375.525 47.76 ;
      RECT 374.525 48.76 375.525 49.76 ;
      RECT 374.525 50.76 375.525 51.76 ;
      RECT 374.525 52.76 375.525 53.76 ;
      RECT 374.525 54.76 375.525 55.76 ;
      RECT 227.52 145.655 228.52 146.655 ;
      RECT 227.52 147.655 228.52 148.655 ;
      RECT 227.52 149.655 228.52 150.655 ;
      RECT 227.52 151.655 228.52 152.655 ;
      RECT 225.52 145.655 226.52 146.655 ;
      RECT 225.52 147.655 226.52 148.655 ;
      RECT 225.52 149.655 226.52 150.655 ;
      RECT 225.52 151.655 226.52 152.655 ;
      RECT 223.52 145.655 224.52 146.655 ;
      RECT 223.52 147.655 224.52 148.655 ;
      RECT 223.52 149.655 224.52 150.655 ;
      RECT 223.52 151.655 224.52 152.655 ;
      RECT 221.52 145.655 222.52 146.655 ;
      RECT 221.52 147.655 222.52 148.655 ;
      RECT 221.52 149.655 222.52 150.655 ;
      RECT 221.52 151.655 222.52 152.655 ;
      RECT 126.925 131.675 127.925 132.675 ;
      RECT 126.925 133.675 127.925 134.675 ;
      RECT 126.925 135.675 127.925 136.675 ;
      RECT 126.925 137.675 127.925 138.675 ;
      RECT 124.925 131.675 125.925 132.675 ;
      RECT 124.925 133.675 125.925 134.675 ;
      RECT 124.925 135.675 125.925 136.675 ;
      RECT 124.925 137.675 125.925 138.675 ;
      RECT 122.925 131.675 123.925 132.675 ;
      RECT 122.925 133.675 123.925 134.675 ;
      RECT 122.925 135.675 123.925 136.675 ;
      RECT 122.925 137.675 123.925 138.675 ;
      RECT 120.925 131.675 121.925 132.675 ;
      RECT 120.925 133.675 121.925 134.675 ;
      RECT 120.925 135.675 121.925 136.675 ;
      RECT 120.925 137.675 121.925 138.675 ;
    LAYER Metal1 ;
      RECT 410.5 46.2 544.75 54.2 ;
      RECT 130.3 31.45 138.3 51.65 ;
      RECT 410.5 31.45 418.5 54.2 ;
      RECT 130.3 31.45 418.5 39.45 ;
      RECT 730 114.765 755 124.765 ;
      RECT 723.165 43.335 749 53.335 ;
      RECT 658.61 131.175 678.425 139.175 ;
      RECT 536.575 199.105 544.575 218.33 ;
      RECT 441.285 22.805 449.285 43.505 ;
      RECT 400 114.765 425 124.765 ;
      RECT 360 46.26 384.025 56.26 ;
      RECT 210.075 145.155 229.02 153.155 ;
      RECT 108.61 131.175 128.425 139.175 ;
  END
END MoS2Xor

MACRO MoS2triNand
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MoS2triNand 0 0 ;
  SIZE 200 BY 280 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 10 0 20 134.05 ;
    END
    PORT
      LAYER NSD ;
        RECT 90 0 100 134.05 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 0 200 20 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Contact ;
        RECT 137.335 216.06 138.335 217.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 137.335 218.06 138.335 219.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 137.335 220.06 138.335 221.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 137.335 222.06 138.335 223.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 137.335 262.115 138.335 263.115 ;
    END
    PORT
      LAYER Contact ;
        RECT 137.335 264.115 138.335 265.115 ;
    END
    PORT
      LAYER Contact ;
        RECT 137.335 266.115 138.335 267.115 ;
    END
    PORT
      LAYER Contact ;
        RECT 137.335 268.115 138.335 269.115 ;
    END
    PORT
      LAYER Contact ;
        RECT 135.335 216.06 136.335 217.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 135.335 218.06 136.335 219.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 135.335 220.06 136.335 221.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 135.335 222.06 136.335 223.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 135.335 262.115 136.335 263.115 ;
    END
    PORT
      LAYER Contact ;
        RECT 135.335 264.115 136.335 265.115 ;
    END
    PORT
      LAYER Contact ;
        RECT 135.335 266.115 136.335 267.115 ;
    END
    PORT
      LAYER Contact ;
        RECT 135.335 268.115 136.335 269.115 ;
    END
    PORT
      LAYER Contact ;
        RECT 133.335 216.06 134.335 217.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 133.335 218.06 134.335 219.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 133.335 220.06 134.335 221.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 133.335 222.06 134.335 223.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 133.335 262.115 134.335 263.115 ;
    END
    PORT
      LAYER Contact ;
        RECT 133.335 264.115 134.335 265.115 ;
    END
    PORT
      LAYER Contact ;
        RECT 133.335 266.115 134.335 267.115 ;
    END
    PORT
      LAYER Contact ;
        RECT 133.335 268.115 134.335 269.115 ;
    END
    PORT
      LAYER Contact ;
        RECT 131.335 216.06 132.335 217.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 131.335 218.06 132.335 219.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 131.335 220.06 132.335 221.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 131.335 222.06 132.335 223.06 ;
    END
    PORT
      LAYER Contact ;
        RECT 131.335 262.115 132.335 263.115 ;
    END
    PORT
      LAYER Contact ;
        RECT 131.335 264.115 132.335 265.115 ;
    END
    PORT
      LAYER Contact ;
        RECT 131.335 266.115 132.335 267.115 ;
    END
    PORT
      LAYER Contact ;
        RECT 131.335 268.115 132.335 269.115 ;
    END
    PORT
      LAYER NSD ;
        RECT 130 170 140 223.58 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 260 200 280 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 130.835 215.56 138.835 269.615 ;
    END
  END VDD
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER NSD ;
        RECT 150 44.03 160 200 ;
    END
  END VOUT
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NSD ;
        RECT 30 170 40 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 70 170 80 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 110 170 120 250 ;
    END
    PORT
      LAYER NSD ;
        RECT 0 230 200 250 ;
    END
  END VSS
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 139 20.55 151 135.05 ;
        RECT 59 20.55 151 32.55 ;
        RECT 59 20.55 71 135.05 ;
    END
  END A
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Gate ;
        RECT 19 139.05 111 149.05 ;
        RECT 99 43.25 111 149.05 ;
        RECT 19 43.45 31 149.05 ;
    END
  END C
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 41.25 35.175 129.165 43.175 ;
      LAYER Gate ;
        RECT 119 43.05 131 135.05 ;
        RECT 121.15 35.2 129.15 135.05 ;
        RECT 39 43.05 51 135.05 ;
        RECT 41.25 35.2 49.25 135.05 ;
      LAYER Cont ;
        RECT 41.75 41.675 42.75 42.675 ;
        RECT 41.75 39.675 42.75 40.675 ;
        RECT 41.75 37.675 42.75 38.675 ;
        RECT 41.75 35.675 42.75 36.675 ;
        RECT 43.75 41.675 44.75 42.675 ;
        RECT 43.75 39.675 44.75 40.675 ;
        RECT 43.75 37.675 44.75 38.675 ;
        RECT 43.75 35.675 44.75 36.675 ;
        RECT 45.75 41.675 46.75 42.675 ;
        RECT 45.75 39.675 46.75 40.675 ;
        RECT 45.75 37.675 46.75 38.675 ;
        RECT 45.75 35.675 46.75 36.675 ;
        RECT 47.75 41.675 48.75 42.675 ;
        RECT 47.75 39.675 48.75 40.675 ;
        RECT 47.75 37.675 48.75 38.675 ;
        RECT 47.75 35.675 48.75 36.675 ;
        RECT 121.665 41.675 122.665 42.675 ;
        RECT 121.665 39.675 122.665 40.675 ;
        RECT 121.665 37.675 122.665 38.675 ;
        RECT 121.665 35.675 122.665 36.675 ;
        RECT 123.665 41.675 124.665 42.675 ;
        RECT 123.665 39.675 124.665 40.675 ;
        RECT 123.665 37.675 124.665 38.675 ;
        RECT 123.665 35.675 124.665 36.675 ;
        RECT 125.665 41.675 126.665 42.675 ;
        RECT 125.665 39.675 126.665 40.675 ;
        RECT 125.665 37.675 126.665 38.675 ;
        RECT 125.665 35.675 126.665 36.675 ;
        RECT 127.665 41.675 128.665 42.675 ;
        RECT 127.665 39.675 128.665 40.675 ;
        RECT 127.665 37.675 128.665 38.675 ;
        RECT 127.665 35.675 128.665 36.675 ;
    END
  END B
  OBS
    LAYER Gate ;
      RECT 79 205 111 215 ;
      RECT 99 155 111 215 ;
      RECT 39 205 71 215 ;
      RECT 59 155 71 215 ;
      RECT 19 155 31 215 ;
      RECT 139 155 151 205.1 ;
      RECT 79 155 91 215 ;
      RECT 39 155 51 215 ;
      RECT 99 155 151 167 ;
      RECT 59 155 91 165 ;
      RECT 19 155 51 165 ;
      RECT 9 206 19 214 ;
      RECT 130 215 139 224 ;
      RECT 130 260 139 270 ;
    LAYER NSD ;
      RECT 10 154.5 20 215.25 ;
      RECT 90 154.5 100 200 ;
      RECT 50 154.5 60 200 ;
      RECT 10 154.5 100 164.5 ;
      RECT 70 44.05 80 164.5 ;
      RECT 130 44.03 140 134.03 ;
      RECT 110 44.03 120 134.03 ;
      RECT 50 44.03 60 134.03 ;
      RECT 30 44.03 40 134.03 ;
      RECT 20 206 29 215 ;
      RECT 41 35 50 44 ;
      RECT 121 35 130 44 ;
    LAYER Contact ;
      RECT 16.555 206.77 17.555 207.77 ;
      RECT 16.555 208.77 17.555 209.77 ;
      RECT 16.555 210.77 17.555 211.77 ;
      RECT 16.555 212.77 17.555 213.77 ;
      RECT 14.555 206.77 15.555 207.77 ;
      RECT 14.555 208.77 15.555 209.77 ;
      RECT 14.555 210.77 15.555 211.77 ;
      RECT 14.555 212.77 15.555 213.77 ;
      RECT 12.555 206.77 13.555 207.77 ;
      RECT 12.555 208.77 13.555 209.77 ;
      RECT 12.555 210.77 13.555 211.77 ;
      RECT 12.555 212.77 13.555 213.77 ;
      RECT 10.555 206.77 11.555 207.77 ;
      RECT 10.555 208.77 11.555 209.77 ;
      RECT 10.555 210.77 11.555 211.77 ;
      RECT 10.555 212.77 11.555 213.77 ;
      RECT 79 205 111 215 ;
      RECT 99 155 111 215 ;
      RECT 39 205 71 215 ;
      RECT 59 155 71 215 ;
      RECT 19 155 31 215 ;
      RECT 139 155 151 205.1 ;
      RECT 79 155 91 215 ;
      RECT 39 155 51 215 ;
      RECT 99 155 151 167 ;
      RECT 59 155 91 165 ;
      RECT 19 155 51 165 ;
        RECT 139 20.55 151 135.05 ;
        RECT 59 20.55 151 32.55 ;
        RECT 59 20.55 71 135.05 ;
        RECT 19 139.05 111 149.05 ;
        RECT 99 43.25 111 149.05 ;
        RECT 19 43.45 31 149.05 ;
        RECT 119 43.05 131 135.05 ;
        RECT 121.15 35.2 129.15 135.05 ;
        RECT 39 43.05 51 135.05 ;
        RECT 41.25 35.2 49.25 135.05 ;
    LAYER Cont ;
      RECT 27.475 206.77 28.475 207.77 ;
      RECT 27.475 208.77 28.475 209.77 ;
      RECT 27.475 210.77 28.475 211.77 ;
      RECT 27.475 212.77 28.475 213.77 ;
      RECT 25.475 206.77 26.475 207.77 ;
      RECT 25.475 208.77 26.475 209.77 ;
      RECT 25.475 210.77 26.475 211.77 ;
      RECT 25.475 212.77 26.475 213.77 ;
      RECT 23.475 206.77 24.475 207.77 ;
      RECT 23.475 208.77 24.475 209.77 ;
      RECT 23.475 210.77 24.475 211.77 ;
      RECT 23.475 212.77 24.475 213.77 ;
      RECT 21.475 206.77 22.475 207.77 ;
      RECT 21.475 208.77 22.475 209.77 ;
      RECT 21.475 210.77 22.475 211.77 ;
      RECT 21.475 212.77 22.475 213.77 ;
      RECT 10 154.5 20 215.25 ;
      RECT 90 154.5 100 200 ;
      RECT 50 154.5 60 200 ;
      RECT 10 154.5 100 164.5 ;
      RECT 70 44.05 80 164.5 ;
      RECT 130 44.03 140 134.03 ;
      RECT 110 44.03 120 134.03 ;
      RECT 50 44.03 60 134.03 ;
      RECT 30 44.03 40 134.03 ;
        RECT 10 0 20 134.05 ;
        RECT 90 0 100 134.05 ;
        RECT 0 0 200 20 ;
        RECT 130 170 140 223.58 ;
        RECT 0 260 200 280 ;
        RECT 150 44.03 160 200 ;
        RECT 30 170 40 250 ;
        RECT 70 170 80 250 ;
        RECT 110 170 120 250 ;
        RECT 0 230 200 250 ;
    LAYER Metal1 ;
      RECT 10.055 206.27 28.975 214.27 ;
  END
END MoS2triNand


END LIBRARY
